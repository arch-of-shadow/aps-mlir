--------------------------------------------------------------------------------
--                  FixRealKCM_Freq200_uid6_T0_Freq200_uid9
-- VHDL generated for DummyFPGA @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq200_uid6_T0_Freq200_uid9 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(19 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq200_uid6_T0_Freq200_uid9 is
signal Y0 :  std_logic_vector(19 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(19 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "00000000000000000010" when "00000",
      "00000110010010001010" when "00001",
      "00001100100100010010" when "00010",
      "00010010110110011010" when "00011",
      "00011001001000100010" when "00100",
      "00011111011010101010" when "00101",
      "00100101101100110010" when "00110",
      "00101011111110111001" when "00111",
      "00110010010001000001" when "01000",
      "00111000100011001001" when "01001",
      "00111110110101010001" when "01010",
      "01000101000111011001" when "01011",
      "01001011011001100001" when "01100",
      "01010001101011101001" when "01101",
      "01010111111101110001" when "01110",
      "01011110001111111001" when "01111",
      "01100100100010000001" when "10000",
      "01101010110100001001" when "10001",
      "01110001000110010001" when "10010",
      "01110111011000011001" when "10011",
      "01111101101010100001" when "10100",
      "10000011111100101000" when "10101",
      "10001010001110110000" when "10110",
      "10010000100000111000" when "10111",
      "10010110110011000000" when "11000",
      "10011101000101001000" when "11001",
      "10100011010111010000" when "11010",
      "10101001101001011000" when "11011",
      "10101111111011100000" when "11100",
      "10110110001101101000" when "11101",
      "10111100011111110000" when "11110",
      "11000010110001111000" when "11111",
      "--------------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                  FixRealKCM_Freq200_uid6_T1_Freq200_uid12
-- VHDL generated for DummyFPGA @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq200_uid6_T1_Freq200_uid12 is
    port (X : in  std_logic_vector(4 downto 0);
          Y : out  std_logic_vector(14 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq200_uid6_T1_Freq200_uid12 is
signal Y0 :  std_logic_vector(14 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(14 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "000000000000000" when "00000",
      "000001100100100" when "00001",
      "000011001001000" when "00010",
      "000100101101101" when "00011",
      "000110010010001" when "00100",
      "000111110110101" when "00101",
      "001001011011001" when "00110",
      "001010111111110" when "00111",
      "001100100100010" when "01000",
      "001110001000110" when "01001",
      "001111101101010" when "01010",
      "010001010001111" when "01011",
      "010010110110011" when "01100",
      "010100011010111" when "01101",
      "010101111111011" when "01110",
      "010111100100000" when "01111",
      "011001001000100" when "10000",
      "011010101101000" when "10001",
      "011100010001100" when "10010",
      "011101110110001" when "10011",
      "011111011010101" when "10100",
      "100000111111001" when "10101",
      "100010100011101" when "10110",
      "100100001000010" when "10111",
      "100101101100110" when "11000",
      "100111010001010" when "11001",
      "101000110101110" when "11010",
      "101010011010011" when "11011",
      "101011111110111" when "11100",
      "101101100011011" when "11101",
      "101111000111111" when "11110",
      "110000101100100" when "11111",
      "---------------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                  FixRealKCM_Freq200_uid6_T2_Freq200_uid15
-- VHDL generated for DummyFPGA @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.600000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq200_uid6_T2_Freq200_uid15 is
    port (X : in  std_logic_vector(5 downto 0);
          Y : out  std_logic_vector(9 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq200_uid6_T2_Freq200_uid15 is
signal Y0 :  std_logic_vector(9 downto 0);
   -- timing of Y0: (c0, 0.600000ns)
signal Y1 :  std_logic_vector(9 downto 0);
   -- timing of Y1: (c0, 0.600000ns)
begin
   with X  select  Y0 <= 
      "0000000000" when "000000",
      "0000001101" when "000001",
      "0000011001" when "000010",
      "0000100110" when "000011",
      "0000110010" when "000100",
      "0000111111" when "000101",
      "0001001011" when "000110",
      "0001011000" when "000111",
      "0001100101" when "001000",
      "0001110001" when "001001",
      "0001111110" when "001010",
      "0010001010" when "001011",
      "0010010111" when "001100",
      "0010100011" when "001101",
      "0010110000" when "001110",
      "0010111100" when "001111",
      "0011001001" when "010000",
      "0011010110" when "010001",
      "0011100010" when "010010",
      "0011101111" when "010011",
      "0011111011" when "010100",
      "0100001000" when "010101",
      "0100010100" when "010110",
      "0100100001" when "010111",
      "0100101110" when "011000",
      "0100111010" when "011001",
      "0101000111" when "011010",
      "0101010011" when "011011",
      "0101100000" when "011100",
      "0101101100" when "011101",
      "0101111001" when "011110",
      "0110000110" when "011111",
      "0110010010" when "100000",
      "0110011111" when "100001",
      "0110101011" when "100010",
      "0110111000" when "100011",
      "0111000100" when "100100",
      "0111010001" when "100101",
      "0111011110" when "100110",
      "0111101010" when "100111",
      "0111110111" when "101000",
      "1000000011" when "101001",
      "1000010000" when "101010",
      "1000011100" when "101011",
      "1000101001" when "101100",
      "1000110101" when "101101",
      "1001000010" when "101110",
      "1001001111" when "101111",
      "1001011011" when "110000",
      "1001101000" when "110001",
      "1001110100" when "110010",
      "1010000001" when "110011",
      "1010001101" when "110100",
      "1010011010" when "110101",
      "1010100111" when "110110",
      "1010110011" when "110111",
      "1011000000" when "111000",
      "1011001100" when "111001",
      "1011011001" when "111010",
      "1011100101" when "111011",
      "1011110010" when "111100",
      "1011111111" when "111101",
      "1100001011" when "111110",
      "1100011000" when "111111",
      "----------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_23_3_Freq200_uid19
-- VHDL generated for DummyFPGA @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X1 X0
-- Output signals: R
--  approx. input signal timings: X1: (c0, 0.000000ns)X0: (c0, 0.000000ns)
--  approx. output signal timings: R: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_23_3_Freq200_uid19 is
    port (X1 : in  std_logic_vector(1 downto 0);
          X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_23_3_Freq200_uid19 is
signal X :  std_logic_vector(4 downto 0);
   -- timing of X: (c0, 0.000000ns)
signal R0 :  std_logic_vector(2 downto 0);
   -- timing of R0: (c0, 0.550000ns)
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100",
      "010" when "00011" | "00101" | "00110" | "01000" | "10000",
      "011" when "00111" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100",
      "100" when "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11000",
      "101" when "01111" | "10111" | "11001" | "11010" | "11100",
      "110" when "11011" | "11101" | "11110",
      "111" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                       Compressor_14_3_Freq200_uid35
-- VHDL generated for DummyFPGA @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X1 X0
-- Output signals: R
--  approx. input signal timings: X1: (c0, 0.000000ns)X0: (c0, 0.000000ns)
--  approx. output signal timings: R: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_14_3_Freq200_uid35 is
    port (X1 : in  std_logic_vector(0 downto 0);
          X0 : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_14_3_Freq200_uid35 is
signal X :  std_logic_vector(4 downto 0);
   -- timing of X: (c0, 0.000000ns)
signal R0 :  std_logic_vector(2 downto 0);
   -- timing of R0: (c0, 0.550000ns)
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10001" | "10010" | "10100" | "11000",
      "100" when "01111" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "101" when "10111" | "11011" | "11101" | "11110",
      "110" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                      FixFunctionByTable_Freq200_uid41
-- Evaluator for x*x on [0,1) for lsbIn=-7 (wIn=7), msbout=-1, lsbOut=-7 (wOut=7). Out interval: [0; 0.984436]. Output is unsigned

-- VHDL generated for DummyFPGA @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2010-2018)
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c0, 0.550000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixFunctionByTable_Freq200_uid41 is
    port (X : in  std_logic_vector(6 downto 0);
          Y : out  std_logic_vector(6 downto 0)   );
end entity;

architecture arch of FixFunctionByTable_Freq200_uid41 is
signal Y0 :  std_logic_vector(6 downto 0);
   -- timing of Y0: (c0, 0.550000ns)
signal Y1 :  std_logic_vector(6 downto 0);
   -- timing of Y1: (c0, 0.550000ns)
begin
   with X  select  Y0 <= 
      "0000000" when "0000000",
      "0000000" when "0000001",
      "0000000" when "0000010",
      "0000000" when "0000011",
      "0000000" when "0000100",
      "0000000" when "0000101",
      "0000000" when "0000110",
      "0000000" when "0000111",
      "0000000" when "0001000",
      "0000001" when "0001001",
      "0000001" when "0001010",
      "0000001" when "0001011",
      "0000001" when "0001100",
      "0000001" when "0001101",
      "0000010" when "0001110",
      "0000010" when "0001111",
      "0000010" when "0010000",
      "0000010" when "0010001",
      "0000011" when "0010010",
      "0000011" when "0010011",
      "0000011" when "0010100",
      "0000011" when "0010101",
      "0000100" when "0010110",
      "0000100" when "0010111",
      "0000100" when "0011000",
      "0000101" when "0011001",
      "0000101" when "0011010",
      "0000110" when "0011011",
      "0000110" when "0011100",
      "0000111" when "0011101",
      "0000111" when "0011110",
      "0001000" when "0011111",
      "0001000" when "0100000",
      "0001001" when "0100001",
      "0001001" when "0100010",
      "0001010" when "0100011",
      "0001010" when "0100100",
      "0001011" when "0100101",
      "0001011" when "0100110",
      "0001100" when "0100111",
      "0001100" when "0101000",
      "0001101" when "0101001",
      "0001110" when "0101010",
      "0001110" when "0101011",
      "0001111" when "0101100",
      "0010000" when "0101101",
      "0010001" when "0101110",
      "0010001" when "0101111",
      "0010010" when "0110000",
      "0010011" when "0110001",
      "0010100" when "0110010",
      "0010100" when "0110011",
      "0010101" when "0110100",
      "0010110" when "0110101",
      "0010111" when "0110110",
      "0011000" when "0110111",
      "0011000" when "0111000",
      "0011001" when "0111001",
      "0011010" when "0111010",
      "0011011" when "0111011",
      "0011100" when "0111100",
      "0011101" when "0111101",
      "0011110" when "0111110",
      "0011111" when "0111111",
      "0100000" when "1000000",
      "0100001" when "1000001",
      "0100010" when "1000010",
      "0100011" when "1000011",
      "0100100" when "1000100",
      "0100101" when "1000101",
      "0100110" when "1000110",
      "0100111" when "1000111",
      "0101000" when "1001000",
      "0101010" when "1001001",
      "0101011" when "1001010",
      "0101100" when "1001011",
      "0101101" when "1001100",
      "0101110" when "1001101",
      "0110000" when "1001110",
      "0110001" when "1001111",
      "0110010" when "1010000",
      "0110011" when "1010001",
      "0110101" when "1010010",
      "0110110" when "1010011",
      "0110111" when "1010100",
      "0111000" when "1010101",
      "0111010" when "1010110",
      "0111011" when "1010111",
      "0111100" when "1011000",
      "0111110" when "1011001",
      "0111111" when "1011010",
      "1000001" when "1011011",
      "1000010" when "1011100",
      "1000100" when "1011101",
      "1000101" when "1011110",
      "1000111" when "1011111",
      "1001000" when "1100000",
      "1001010" when "1100001",
      "1001011" when "1100010",
      "1001101" when "1100011",
      "1001110" when "1100100",
      "1010000" when "1100101",
      "1010001" when "1100110",
      "1010011" when "1100111",
      "1010100" when "1101000",
      "1010110" when "1101001",
      "1011000" when "1101010",
      "1011001" when "1101011",
      "1011011" when "1101100",
      "1011101" when "1101101",
      "1011111" when "1101110",
      "1100000" when "1101111",
      "1100010" when "1110000",
      "1100100" when "1110001",
      "1100110" when "1110010",
      "1100111" when "1110011",
      "1101001" when "1110100",
      "1101011" when "1110101",
      "1101101" when "1110110",
      "1101111" when "1110111",
      "1110000" when "1111000",
      "1110010" when "1111001",
      "1110100" when "1111010",
      "1110110" when "1111011",
      "1111000" when "1111100",
      "1111010" when "1111101",
      "1111100" when "1111110",
      "1111110" when "1111111",
      "-------" when others;
   Y1 <= Y0; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                          SinCosTable_Freq200_uid4
-- VHDL generated for DummyFPGA @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.550000ns)
--  approx. output signal timings: Y: (c1, 2.789062ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity SinCosTable_Freq200_uid4 is
    port (clk, rst : in std_logic;
          X : in  std_logic_vector(9 downto 0);
          Y : out  std_logic_vector(55 downto 0)   );
end entity;

architecture arch of SinCosTable_Freq200_uid4 is
signal Y0, Y0_d1 :  std_logic_vector(55 downto 0);
   -- timing of Y0: (c0, 2.550000ns)
signal Y1 :  std_logic_vector(55 downto 0);
   -- timing of Y1: (c1, 2.789062ns)
begin
   process(clk, rst)
      begin
         if rst = '1' then
            Y0_d1 <=  (others => '0');
         elsif clk'event and clk = '1' then
            Y0_d1 <=  Y0;
         end if;
      end process;
   with X  select  Y0 <= 
      "00000000000000000000000010001111111111111111111111111000" when "0000000000",
      "00000000001100100100010001111111111111111111111110101001" when "0000000001",
      "00000000011001001000100001111111111111111111111010111100" when "0000000010",
      "00000000100101101100110001101111111111111111110100110001" when "0000000011",
      "00000000110010010001000001001111111111111111101100001001" when "0000000100",
      "00000000111110110101010000101111111111111111100001000010" when "0000000101",
      "00000001001011011001100000001111111111111111010011011110" when "0000000110",
      "00000001010111111101101111011111111111111111000011011011" when "0000000111",
      "00000001100100100001111110011111111111111110110000111011" when "0000001000",
      "00000001110001000110001101001111111111111110011011111101" when "0000001001",
      "00000001111101101010011011101111111111111110000100100000" when "0000001010",
      "00000010001010001110101001111111111111111101101010100110" when "0000001011",
      "00000010010110110010110111101111111111111101001110001110" when "0000001100",
      "00000010100011010111000101001111111111111100101111011000" when "0000001101",
      "00000010101111111011010010001111111111111100001110000101" when "0000001110",
      "00000010111100011111011110111111111111111011101010010011" when "0000001111",
      "00000011001001000011101011001111111111111011000100000011" when "0000010000",
      "00000011010101100111110110111111111111111010011011010110" when "0000010001",
      "00000011100010001100000010001111111111111001110000001010" when "0000010010",
      "00000011101110110000001100101111111111111001000010100001" when "0000010011",
      "00000011111011010100010110111111111111111000010010011010" when "0000010100",
      "00000100000111111000100000011111111111110111011111110101" when "0000010101",
      "00000100010100011100101001001111111111110110101010110010" when "0000010110",
      "00000100100001000000110001011111111111110101110011010001" when "0000010111",
      "00000100101101100100111000111111111111110100111001010010" when "0000011000",
      "00000100111010001000111111101111111111110011111100110101" when "0000011001",
      "00000101000110101101000101101111111111110010111101111011" when "0000011010",
      "00000101010011010001001010111111111111110001111100100011" when "0000011011",
      "00000101011111110101001111001111111111110000111000101100" when "0000011100",
      "00000101101100011001010010101111111111101111110010011000" when "0000011101",
      "00000101111000111101010101011111111111101110101001100110" when "0000011110",
      "00000110000101100001010111001111111111101101011110010110" when "0000011111",
      "00000110010010000101010111111111111111101100010000101000" when "0000100000",
      "00000110011110101001010111111111111111101011000000011101" when "0000100001",
      "00000110101011001101010110101111111111101001101101110011" when "0000100010",
      "00000110110111110001010100101111111111101000011000101100" when "0000100011",
      "00000111000100010101010001011111111111100111000001000110" when "0000100100",
      "00000111010000111001001100111111111111100101100111000011" when "0000100101",
      "00000111011101011101000111101111111111100100001010100010" when "0000100110",
      "00000111101010000001000000111111111111100010101011100100" when "0000100111",
      "00000111110110100100111001001111111111100001001010000111" when "0000101000",
      "00001000000011001000110000001111111111011111100110001101" when "0000101001",
      "00001000001111101100100101111111111111011101111111110100" when "0000101010",
      "00001000011100010000011010011111111111011100010110111110" when "0000101011",
      "00001000101000110100001101101111111111011010101011101010" when "0000101100",
      "00001000110101010111111111101111111111011000111101111000" when "0000101101",
      "00001001000001111011110000001111111111010111001101101001" when "0000101110",
      "00001001001110011111011111001111111111010101011010111011" when "0000101111",
      "00001001011011000011001100111111111111010011100101110000" when "0000110000",
      "00001001100111100110111001001111111111010001101110000111" when "0000110001",
      "00001001110100001010100011111111111111001111110100000000" when "0000110010",
      "00001010000000101110001101001111111111001101110111011011" when "0000110011",
      "00001010001101010001110100111111111111001011111000011001" when "0000110100",
      "00001010011001110101011010111111111111001001110110111001" when "0000110101",
      "00001010100110011000111111011111111111000111110010111011" when "0000110110",
      "00001010110010111100100010011111111111000101101100011111" when "0000110111",
      "00001010111111100000000011101111111111000011100011100101" when "0000111000",
      "00001011001100000011100011001111111111000001011000001110" when "0000111001",
      "00001011011000100111000000111111111110111111001010011001" when "0000111010",
      "00001011100101001010011100111111111110111100111010000110" when "0000111011",
      "00001011110001101101110111001111111110111010100111010110" when "0000111100",
      "00001011111110010001001111101111111110111000010010000111" when "0000111101",
      "00001100001010110100100110011111111110110101111010011011" when "0000111110",
      "00001100010111010111111010111111111110110011100000010001" when "0000111111",
      "00001100100011111011001101111111111110110001000011101010" when "0001000000",
      "00001100110000011110011110101111111110101110100100100100" when "0001000001",
      "00001100111101000001101101101111111110101100000011000001" when "0001000010",
      "00001101001001100100111010101111111110101001011111000001" when "0001000011",
      "00001101010110001000000101011111111110100110111000100010" when "0001000100",
      "00001101100010101011001110001111111110100100001111100110" when "0001000101",
      "00001101101111001110010100111111111110100001100100001100" when "0001000110",
      "00001101111011110001011001101111111110011110110110010101" when "0001000111",
      "00001110001000010100011100001111111110011100000110000000" when "0001001000",
      "00001110010100110111011100011111111110011001010011001101" when "0001001001",
      "00001110100001011010011010011111111110010110011101111100" when "0001001010",
      "00001110101101111101010110011111111110010011100110001110" when "0001001011",
      "00001110111010100000001111111111111110010000101100000010" when "0001001100",
      "00001111000111000011000111001111111110001101101111011001" when "0001001101",
      "00001111010011100101111100001111111110001010110000010010" when "0001001110",
      "00001111100000001000101110101111111110000111101110101101" when "0001001111",
      "00001111101100101011011110111111111110000100101010101011" when "0001010000",
      "00001111111001001110001100101111111110000001100100001011" when "0001010001",
      "00010000000101110000110111111111111101111110011011001101" when "0001010010",
      "00010000010010010011100000111111111101111011001111110010" when "0001010011",
      "00010000011110110110000111001111111101111000000001111001" when "0001010100",
      "00010000101011011000101010111111111101110100110001100011" when "0001010101",
      "00010000110111111011001100001111111101110001011110101111" when "0001010110",
      "00010001000100011101101010101111111101101110001001011101" when "0001010111",
      "00010001010001000000000110101111111101101010110001101110" when "0001011000",
      "00010001011101100010011111111111111101100111010111100010" when "0001011001",
      "00010001101010000100110110101111111101100011111010111000" when "0001011010",
      "00010001110110100111001010101111111101100000011011110000" when "0001011011",
      "00010010000011001001011011101111111101011100111010001011" when "0001011100",
      "00010010001111101011101010001111111101011001010110001000" when "0001011101",
      "00010010011100001101110101101111111101010101101111101000" when "0001011110",
      "00010010101000101111111110011111111101010010000110101010" when "0001011111",
      "00010010110101010010000100001111111101001110011011001111" when "0001100000",
      "00010011000001110100000111001111111101001010101101010110" when "0001100001",
      "00010011001110010110000111001111111101000110111101000000" when "0001100010",
      "00010011011010111000000100001111111101000011001010001100" when "0001100011",
      "00010011100111011001111110001111111100111111010100111011" when "0001100100",
      "00010011110011111011110101001111111100111011011101001100" when "0001100101",
      "00010100000000011101101001001111111100110111100011000000" when "0001100110",
      "00010100001100111111011001111111111100110011100110010111" when "0001100111",
      "00010100011001100001000111101111111100101111100111010000" when "0001101000",
      "00010100100110000010110010011111111100101011100101101011" when "0001101001",
      "00010100110010100100011001101111111100100111100001101010" when "0001101010",
      "00010100111111000101111101111111111100100011011011001011" when "0001101011",
      "00010101001011100111011110111111111100011111010010001110" when "0001101100",
      "00010101011000001000111100101111111100011011000110110100" when "0001101101",
      "00010101100100101010010111001111111100010110111000111101" when "0001101110",
      "00010101110001001011101110001111111100010010101000101000" when "0001101111",
      "00010101111101101101000001111111111100001110010101110110" when "0001110000",
      "00010110001010001110010010011111111100001010000000100111" when "0001110001",
      "00010110010110101111011111001111111100000101101000111011" when "0001110010",
      "00010110100011010000101000101111111100000001001110110001" when "0001110011",
      "00010110101111110001101110101111111011111100110010001010" when "0001110100",
      "00010110111100010010110001011111111011111000010011000101" when "0001110101",
      "00010111001000110011110000001111111011110011110001100011" when "0001110110",
      "00010111010101010100101011101111111011101111001101100100" when "0001110111",
      "00010111100001110101100011011111111011101010100111001000" when "0001111000",
      "00010111101110010110010111101111111011100101111110001111" when "0001111001",
      "00010111111010110111001000001111111011100001010010111000" when "0001111010",
      "00011000000111010111110100111111111011011100100101000100" when "0001111011",
      "00011000010011111000011110001111111011010111110100110011" when "0001111100",
      "00011000100000011001000011011111111011010011000010000100" when "0001111101",
      "00011000101100111001100100111111111011001110001100111001" when "0001111110",
      "00011000111001011010000010101111111011001001010101010000" when "0001111111",
      "00011001000101111010011100101111111011000100011011001010" when "0010000000",
      "00011001010010011010110010101111111010111111011110100111" when "0010000001",
      "00011001011110111011000100111111111010111010011111100111" when "0010000010",
      "00011001101011011011010011001111111010110101011110001001" when "0010000011",
      "00011001110111111011011101011111111010110000011010001111" when "0010000100",
      "00011010000100011011100011101111111010101011010011110111" when "0010000101",
      "00011010010000111011100101111111111010100110001011000011" when "0010000110",
      "00011010011101011011100100001111111010100000111111110001" when "0010000111",
      "00011010101001111011011110011111111010011011110010000010" when "0010001000",
      "00011010110110011011010100011111111010010110100001110110" when "0010001001",
      "00011011000010111011000110001111111010010001001111001101" when "0010001010",
      "00011011001111011010110011111111111010001011111010000111" when "0010001011",
      "00011011011011111010011101011111111010000110100010100101" when "0010001100",
      "00011011101000011010000010101111111010000001001000100101" when "0010001101",
      "00011011110100111001100011101111111001111011101100001000" when "0010001110",
      "00011100000001011001000000011111111001110110001101001110" when "0010001111",
      "00011100001101111000011000111111111001110000101011110111" when "0010010000",
      "00011100011010010111101100111111111001101011001000000011" when "0010010001",
      "00011100100110110110111100101111111001100101100001110010" when "0010010010",
      "00011100110011010110000111111111111001011111111001000100" when "0010010011",
      "00011100111111110101001110101111111001011010001101111010" when "0010010100",
      "00011101001100010100010000111111111001010100100000010010" when "0010010101",
      "00011101011000110011001110111111111001001110110000001110" when "0010010110",
      "00011101100101010010001000001111111001001000111101101101" when "0010010111",
      "00011101110001110000111100111111111001000011001000101111" when "0010011000",
      "00011101111110001111101100111111111000111101010001010100" when "0010011001",
      "00011110001010101110011000101111111000110111010111011100" when "0010011010",
      "00011110010111001100111111011111111000110001011011000111" when "0010011011",
      "00011110100011101011100001101111111000101011011100010110" when "0010011100",
      "00011110110000001001111111001111111000100101011011001000" when "0010011101",
      "00011110111100101000010111111111111000011111010111011101" when "0010011110",
      "00011111001001000110101011111111111000011001010001010101" when "0010011111",
      "00011111010101100100111010111111111000010011001000110001" when "0010100000",
      "00011111100010000011000101011111111000001100111101101111" when "0010100001",
      "00011111101110100001001010111111111000000110110000010001" when "0010100010",
      "00011111111010111111001011011111111000000000100000010111" when "0010100011",
      "00100000000111011101000111001111110111111010001110000000" when "0010100100",
      "00100000010011111010111101101111110111110011111001001100" when "0010100101",
      "00100000100000011000101111011111110111101101100001111011" when "0010100110",
      "00100000101100110110011100001111110111100111001000001110" when "0010100111",
      "00100000111001010100000011111111110111100000101100000100" when "0010101000",
      "00100001000101110001100110011111110111011010001101011110" when "0010101001",
      "00100001010010001111000011111111110111010011101100011011" when "0010101010",
      "00100001011110101100011100011111110111001101001000111011" when "0010101011",
      "00100001101011001001101111011111110111000110100010111111" when "0010101100",
      "00100001110111100110111101011111110110111111111010100110" when "0010101101",
      "00100010000100000100000110011111110110111001001111110001" when "0010101110",
      "00100010010000100001001001111111110110110010100010011111" when "0010101111",
      "00100010011100111110001000001111110110101011110010110001" when "0010110000",
      "00100010101001011011000000111111110110100101000000100110" when "0010110001",
      "00100010110101110111110100101111110110011110001011111111" when "0010110010",
      "00100011000010010100100010111111110110010111010100111011" when "0010110011",
      "00100011001110110001001011101111110110010000011011011011" when "0010110100",
      "00100011011011001101101110111111110110001001011111011111" when "0010110101",
      "00100011100111101010001100111111110110000010100001000110" when "0010110110",
      "00100011110100000110100101011111110101111011100000010001" when "0010110111",
      "00100100000000100010111000001111110101110100011100111111" when "0010111000",
      "00100100001100111111000101101111110101101101010111010001" when "0010111001",
      "00100100011001011011001101011111110101100110001111000111" when "0010111010",
      "00100100100101110111001111011111110101011111000100100001" when "0010111011",
      "00100100110010010011001011111111110101010111110111011110" when "0010111100",
      "00100100111110101111000010111111110101010000100111111111" when "0010111101",
      "00100101001011001010110011111111110101001001010110000011" when "0010111110",
      "00100101010111100110011111011111110101000010000001101100" when "0010111111",
      "00100101100100000010000100111111110100111010101010111000" when "0011000000",
      "00100101110000011101100100111111110100110011010001101000" when "0011000001",
      "00100101111100111000111110111111110100101011110101111011" when "0011000010",
      "00100110001001010100010011001111110100100100010111110011" when "0011000011",
      "00100110010101101111100001011111110100011100110111001110" when "0011000100",
      "00100110100010001010101001101111110100010101010100001110" when "0011000101",
      "00100110101110100101101100001111110100001101101110110001" when "0011000110",
      "00100110111011000000101000101111110100000110000110111000" when "0011000111",
      "00100111000111011011011111001111110011111110011100100011" when "0011001000",
      "00100111010011110110001111011111110011110110101111110010" when "0011001001",
      "00100111100000010000111001111111110011101111000000100101" when "0011001010",
      "00100111101100101011011110001111110011100111001110111100" when "0011001011",
      "00100111111001000101111100001111110011011111011010110111" when "0011001100",
      "00101000000101100000010100001111110011010111100100010110" when "0011001101",
      "00101000010001111010100110001111110011001111101011011001" when "0011001110",
      "00101000011110010100110001101111110011000111110000000000" when "0011001111",
      "00101000101010101110110111001111110010111111110010001011" when "0011010000",
      "00101000110111001000110110001111110010110111110001111010" when "0011010001",
      "00101001000011100010101110111111110010101111101111001101" when "0011010010",
      "00101001001111111100100001011111110010100111101010000100" when "0011010011",
      "00101001011100010110001101011111110010011111100010100000" when "0011010100",
      "00101001101000101111110011001111110010010111011000100000" when "0011010101",
      "00101001110101001001010010011111110010001111001100000100" when "0011010110",
      "00101010000001100010101011011111110010000110111101001100" when "0011010111",
      "00101010001101111011111101101111110001111110101011111000" when "0011011000",
      "00101010011010010101001001011111110001110110011000001001" when "0011011001",
      "00101010100110101110001110111111110001101110000001111110" when "0011011010",
      "00101010110011000111001101101111110001100101101001010111" when "0011011011",
      "00101010111111100000000101101111110001011101001110010100" when "0011011100",
      "00101011001011111000110111001111110001010100110000110110" when "0011011101",
      "00101011011000010001100001111111110001001100010000111100" when "0011011110",
      "00101011100100101010000110001111110001000011101110100111" when "0011011111",
      "00101011110001000010100011101111110000111011001001110101" when "0011100000",
      "00101011111101011010111010011111110000110010100010101001" when "0011100001",
      "00101100001001110011001010001111110000101001111001000001" when "0011100010",
      "00101100010110001011010011011111110000100001001100111101" when "0011100011",
      "00101100100010100011010101101111110000011000011110011101" when "0011100100",
      "00101100101110111011010000111111110000001111101101100011" when "0011100101",
      "00101100111011010011000101011111110000000110111010001100" when "0011100110",
      "00101101000111101010110010111111101111111110000100011010" when "0011100111",
      "00101101010100000010011001101111101111110101001100001101" when "0011101000",
      "00101101100000011001111001001111101111101100010001100101" when "0011101001",
      "00101101101100110001010001111111101111100011010100100001" when "0011101010",
      "00101101111001001000100011011111101111011010010101000001" when "0011101011",
      "00101110000101011111101101111111101111010001010011000110" when "0011101100",
      "00101110010001110110110001001111101111001000001110110000" when "0011101101",
      "00101110011110001101101101011111101110111111000111111111" when "0011101110",
      "00101110101010100100100010011111101110110101111110110010" when "0011101111",
      "00101110110110111011010000011111101110101100110011001010" when "0011110000",
      "00101111000011010001110110111111101110100011100101000111" when "0011110001",
      "00101111001111101000010110011111101110011010010100101000" when "0011110010",
      "00101111011011111110101110011111101110010001000001101111" when "0011110011",
      "00101111101000010100111111011111101110000111101100011010" when "0011110100",
      "00101111110100101011001000101111101101111110010100101010" when "0011110101",
      "00110000000001000001001010111111101101110100111010011111" when "0011110110",
      "00110000001101010111000101011111101101101011011101111001" when "0011110111",
      "00110000011001101100111000101111101101100001111110110111" when "0011111000",
      "00110000100110000010100100011111101101011000011101011011" when "0011111001",
      "00110000110010011000001000101111101101001110111001100011" when "0011111010",
      "00110000111110101101100101011111101101000101010011010001" when "0011111011",
      "00110001001011000010111010101111101100111011101010100100" when "0011111100",
      "00110001010111011000001000001111101100110001111111011011" when "0011111101",
      "00110001100011101101001110001111101100101000010001111000" when "0011111110",
      "00110001110000000010001100101111101100011110100001111001" when "0011111111",
      "00110001111100010111000011001111101100010100101111100000" when "0100000000",
      "00110010001000101011110010001111101100001010111010101100" when "0100000001",
      "00110010010101000000011001011111101100000001000011011101" when "0100000010",
      "00110010100001010100111000111111101011110111001001110100" when "0100000011",
      "00110010101101101001010000101111101011101101001101101111" when "0100000100",
      "00110010111001111101100000101111101011100011001111010000" when "0100000101",
      "00110011000110010001101000101111101011011001001110010101" when "0100000110",
      "00110011010010100101101000101111101011001111001011000001" when "0100000111",
      "00110011011110111001100000111111101011000101000101010001" when "0100001000",
      "00110011101011001101010001001111101010111010111101000111" when "0100001001",
      "00110011110111100000111001101111101010110000110010100010" when "0100001010",
      "00110100000011110100011001111111101010100110100101100010" when "0100001011",
      "00110100010000000111110010001111101010011100010110001000" when "0100001100",
      "00110100011100011011000010011111101010010010000100010011" when "0100001101",
      "00110100101000101110001010101111101010000111110000000100" when "0100001110",
      "00110100110101000001001010101111101001111101011001011010" when "0100001111",
      "00110101000001010100000010011111101001110011000000010110" when "0100010000",
      "00110101001101100110110010001111101001101000100100110111" when "0100010001",
      "00110101011001111001011001101111101001011110000110111110" when "0100010010",
      "00110101100110001011111000111111101001010011100110101010" when "0100010011",
      "00110101110010011110001111111111101001001001000011111100" when "0100010100",
      "00110101111110110000011110101111101000111110011110110011" when "0100010101",
      "00110110001011000010100101001111101000110011110111010000" when "0100010110",
      "00110110010111010100100011001111101000101001001101010011" when "0100010111",
      "00110110100011100110011000101111101000011110100000111011" when "0100011000",
      "00110110101111111000000101111111101000010011110010001001" when "0100011001",
      "00110110111100001001101010111111101000001001000000111101" when "0100011010",
      "00110111001000011011000111001111100111111110001101010111" when "0100011011",
      "00110111010100101100011010111111100111110011010111010110" when "0100011100",
      "00110111100000111101100110001111100111101000011110111100" when "0100011101",
      "00110111101101001110101000111111100111011101100100000111" when "0100011110",
      "00110111111001011111100011001111100111010010100110111000" when "0100011111",
      "00111000000101110000010100101111100111000111100111001111" when "0100100000",
      "00111000010010000000111101011111100110111100100101001011" when "0100100001",
      "00111000011110010001011101101111100110110001100000101110" when "0100100010",
      "00111000101010100001110101001111100110100110011001110111" when "0100100011",
      "00111000110110110010000011111111100110011011010000100110" when "0100100100",
      "00111001000011000010001001111111100110010000000100111010" when "0100100101",
      "00111001001111010010000110111111100110000100110110110101" when "0100100110",
      "00111001011011100001111011011111100101111001100110010110" when "0100100111",
      "00111001100111110001100110111111100101101110010011011101" when "0100101000",
      "00111001110100000001001001011111100101100010111110001010" when "0100101001",
      "00111010000000010000100011001111100101010111100110011101" when "0100101010",
      "00111010001100011111110011111111100101001100001100010111" when "0100101011",
      "00111010011000101110111011101111100101000000101111110111" when "0100101100",
      "00111010100100111101111010011111100100110101010000111101" when "0100101101",
      "00111010110001001100110000001111100100101001101111101001" when "0100101110",
      "00111010111101011011011100111111100100011110001011111011" when "0100101111",
      "00111011001001101010000000011111100100010010100101110100" when "0100110000",
      "00111011010101111000011010111111100100000110111101010011" when "0100110001",
      "00111011100010000110101100001111100011111011010010011001" when "0100110010",
      "00111011101110010100110100001111100011101111100101000101" when "0100110011",
      "00111011111010100010110011001111100011100011110101011000" when "0100110100",
      "00111100000110110000101000111111100011011000000011010000" when "0100110101",
      "00111100010010111110010101001111100011001100001110110000" when "0100110110",
      "00111100011111001011111000011111100011000000010111110110" when "0100110111",
      "00111100101011011001010010001111100010110100011110100010" when "0100111000",
      "00111100110111100110100010101111100010101000100010110110" when "0100111001",
      "00111101000011110011101001101111100010011100100100101111" when "0100111010",
      "00111101010000000000100111001111100010010000100100010000" when "0100111011",
      "00111101011100001101011011011111100010000100100001010111" when "0100111100",
      "00111101101000011010000110001111100001111000011100000100" when "0100111101",
      "00111101110100100110100111001111100001101100010100011001" when "0100111110",
      "00111110000000110010111110111111100001100000001010010100" when "0100111111",
      "00111110001100111111001101001111100001010011111101110110" when "0101000000",
      "00111110011001001011010001101111100001000111101110111111" when "0101000001",
      "00111110100101010111001100011111100000111011011101101111" when "0101000010",
      "00111110110001100010111101101111100000101111001010000101" when "0101000011",
      "00111110111101101110100101001111100000100010110100000011" when "0101000100",
      "00111111001001111010000011001111100000010110011011100111" when "0101000101",
      "00111111010110000101010111001111100000001010000000110011" when "0101000110",
      "00111111100010010000100001011111011111111101100011100101" when "0101000111",
      "00111111101110011011100001111111011111110001000011111111" when "0101001000",
      "00111111111010100110011000101111011111100100100001111111" when "0101001001",
      "01000000000110110001000101101111011111010111111101100111" when "0101001010",
      "01000000010010111011101000011111011111001011010110110101" when "0101001011",
      "01000000011111000110000001101111011110111110101101101011" when "0101001100",
      "01000000101011010000010000101111011110110010000010001000" when "0101001101",
      "01000000110111011010010101111111011110100101010100001100" when "0101001110",
      "01000001000011100100010000111111011110011000100011111000" when "0101001111",
      "01000001001111101110000001111111011110001011110001001010" when "0101010000",
      "01000001011011110111101001001111011101111110111100000101" when "0101010001",
      "01000001101000000001000101111111011101110010000100100110" when "0101010010",
      "01000001110100001010011000111111011101100101001010101111" when "0101010011",
      "01000010000000010011100001011111011101011000001110011111" when "0101010100",
      "01000010001100011100011111111111011101001011001111110110" when "0101010101",
      "01000010011000100101010100001111011100111110001110110101" when "0101010110",
      "01000010100100101101111110011111011100110001001011011100" when "0101010111",
      "01000010110000110110011110001111011100100100000101101010" when "0101011000",
      "01000010111100111110110011101111011100010110111101011111" when "0101011001",
      "01000011001001000110111110101111011100001001110010111100" when "0101011010",
      "01000011010101001110111111101111011011111100100110000001" when "0101011011",
      "01000011100001010110110101111111011011101111010110101110" when "0101011100",
      "01000011101101011110100001111111011011100010000101000010" when "0101011101",
      "01000011111001100110000011101111011011010100110000111101" when "0101011110",
      "01000100000101101101011010101111011011000111011010100001" when "0101011111",
      "01000100010001110100100111001111011010111010000001101100" when "0101100000",
      "01000100011101111011101001011111011010101100100110011111" when "0101100001",
      "01000100101010000010100000111111011010011111001000111010" when "0101100010",
      "01000100110110001001001101101111011010010001101000111101" when "0101100011",
      "01000101000010001111110000001111011010000100000110101000" when "0101100100",
      "01000101001110010110000111101111011001110110100001111011" when "0101100101",
      "01000101011010011100010100101111011001101000111010110101" when "0101100110",
      "01000101100110100010010110111111011001011011010001011000" when "0101100111",
      "01000101110010101000001110101111011001001101100101100010" when "0101101000",
      "01000101111110101101111011011111011000111111110111010101" when "0101101001",
      "01000110001010110011011101011111011000110010000110110000" when "0101101010",
      "01000110010110111000110100011111011000100100010011110011" when "0101101011",
      "01000110100010111110000000111111011000010110011110011110" when "0101101100",
      "01000110101111000011000010001111011000001000100110110010" when "0101101101",
      "01000110111011000111111000101111010111111010101100101101" when "0101101110",
      "01000111000111001100100100011111010111101100110000010001" when "0101101111",
      "01000111010011010001000100111111010111011110110001011101" when "0101110000",
      "01000111011111010101011010101111010111010000110000010010" when "0101110001",
      "01000111101011011001100101001111010111000010101100101110" when "0101110010",
      "01000111110111011101100100111111010110110100100110110100" when "0101110011",
      "01001000000011100001011001001111010110100110011110100001" when "0101110100",
      "01001000001111100101000010101111010110011000010011110111" when "0101110101",
      "01001000011011101000100000111111010110001010000110110110" when "0101110110",
      "01001000100111101011110011111111010101111011110111011101" when "0101110111",
      "01001000110011101110111011101111010101101101100101101101" when "0101111000",
      "01001000111111110001111000011111010101011111010001100101" when "0101111001",
      "01001001001011110100101001101111010101010000111011000111" when "0101111010",
      "01001001010111110111001111111111010101000010100010010000" when "0101111011",
      "01001001100011111001101010101111010100110100000111000011" when "0101111100",
      "01001001101111111011111001111111010100100101101001011110" when "0101111101",
      "01001001111011111101111110001111010100010111001001100010" when "0101111110",
      "01001010000111111111110110101111010100001000100111001110" when "0101111111",
      "01001010010100000001100011111111010011111010000010100100" when "0110000000",
      "01001010100000000011000101101111010011101011011011100011" when "0110000001",
      "01001010101100000100011011111111010011011100110010001010" when "0110000010",
      "01001010111000000101100110101111010011001110000110011010" when "0110000011",
      "01001011000100000110100101111111010010111111011000010100" when "0110000100",
      "01001011010000000111011001011111010010110000100111110110" when "0110000101",
      "01001011011100001000000001101111010010100001110101000010" when "0110000110",
      "01001011101000001000011101111111010010010010111111110110" when "0110000111",
      "01001011110100001000101110101111010010000100001000010100" when "0110001000",
      "01001100000000001000110011101111010001110101001110011011" when "0110001001",
      "01001100001100001000101100111111010001100110010010001011" when "0110001010",
      "01001100011000001000011010101111010001010111010011100100" when "0110001011",
      "01001100100100000111111100011111010001001000010010100111" when "0110001100",
      "01001100110000000111010010011111010000111001001111010010" when "0110001101",
      "01001100111100000110011100011111010000101010001001101000" when "0110001110",
      "01001101001000000101011010101111010000011011000001100110" when "0110001111",
      "01001101010100000100001101001111010000001011110111001110" when "0110010000",
      "01001101100000000010110011101111001111111100101010100000" when "0110010001",
      "01001101101100000001001110001111001111101101011011011011" when "0110010010",
      "01001101110111111111011100101111001111011110001001111111" when "0110010011",
      "01001110000011111101011111001111001111001110110110001110" when "0110010100",
      "01001110001111111011010101101111001110111111100000000101" when "0110010101",
      "01001110011011111001000000001111001110110000000111100111" when "0110010110",
      "01001110100111110110011110011111001110100000101100110010" when "0110010111",
      "01001110110011110011110000101111001110010001001111100110" when "0110011000",
      "01001110111111110000110110101111001110000001110000000101" when "0110011001",
      "01001111001011101101110000011111001101110010001110001101" when "0110011010",
      "01001111010111101010011110001111001101100010101001111111" when "0110011011",
      "01001111100011100110111111011111001101010011000011011011" when "0110011100",
      "01001111101111100011010100101111001101000011011010100001" when "0110011101",
      "01001111111011011111011101011111001100110011101111010001" when "0110011110",
      "01010000000111011011011001111111001100100100000001101011" when "0110011111",
      "01010000010011010111001010001111001100010100010001101111" when "0110100000",
      "01010000011111010010101101111111001100000100011111011101" when "0110100001",
      "01010000101011001110000101011111001011110100101010110101" when "0110100010",
      "01010000110111001001010000001111001011100100110011110111" when "0110100011",
      "01010001000011000100001110101111001011010100111010100011" when "0110100100",
      "01010001001110111111000000101111001011000100111110111010" when "0110100101",
      "01010001011010111001100110001111001010110101000000111011" when "0110100110",
      "01010001100110110011111110111111001010100101000000100110" when "0110100111",
      "01010001110010101110001011001111001010010100111101111011" when "0110101000",
      "01010001111110101000001010111111001010000100111000111011" when "0110101001",
      "01010010001010100001111101111111001001110100110001100101" when "0110101010",
      "01010010010110011011100100001111001001100100100111111010" when "0110101011",
      "01010010100010010100111101111111001001010100011011111001" when "0110101100",
      "01010010101110001110001010111111001001000100001101100010" when "0110101101",
      "01010010111010000111001011001111001000110011111100110110" when "0110101110",
      "01010011000101111111111110011111001000100011101001110101" when "0110101111",
      "01010011010001111000100100111111001000010011010100011110" when "0110110000",
      "01010011011101110000111110101111001000000010111100110011" when "0110110001",
      "01010011101001101001001011101111000111110010100010110001" when "0110110010",
      "01010011110101100001001011101111000111100010000110011011" when "0110110011",
      "01010100000001011000111110101111000111010001100111101111" when "0110110100",
      "01010100001101010000100100101111000111000001000110101110" when "0110110101",
      "01010100011001000111111101101111000110110000100011011000" when "0110110110",
      "01010100100100111111001001111111000110011111111101101101" when "0110110111",
      "01010100110000110110001000111111000110001111010101101101" when "0110111000",
      "01010100111100101100111010111111000101111110101011011000" when "0110111001",
      "01010101001000100011011111101111000101101101111110101110" when "0110111010",
      "01010101010100011001110111011111000101011101001111101111" when "0110111011",
      "01010101100000010000000001111111000101001100011110011011" when "0110111100",
      "01010101101100000101111111011111000100111011101010110010" when "0110111101",
      "01010101110111111011101111101111000100101010110100110101" when "0110111110",
      "01010110000011110001010010011111000100011001111100100010" when "0110111111",
      "01010110001111100110101000001111000100001001000001111011" when "0111000000",
      "01010110011011011011110000011111000011111000000101000000" when "0111000001",
      "01010110100111010000101011101111000011100111000101101111" when "0111000010",
      "01010110110011000101011001001111000011010110000100001010" when "0111000011",
      "01010110111110111001111001011111000011000101000000010001" when "0111000100",
      "01010111001010101110001100011111000010110011111010000011" when "0111000101",
      "01010111010110100010010001111111000010100010110001100000" when "0111000110",
      "01010111100010010110001001111111000010010001100110101001" when "0111000111",
      "01010111101110001001110100001111000010000000011001011110" when "0111001000",
      "01010111111001111101010001001111000001101111001001111110" when "0111001001",
      "01011000000101110000100000101111000001011101111000001010" when "0111001010",
      "01011000010001100011100010011111000001001100100100000010" when "0111001011",
      "01011000011101010110010110101111000000111011001101100110" when "0111001100",
      "01011000101001001000111101001111000000101001110100110101" when "0111001101",
      "01011000110100111011010101111111000000011000011001110000" when "0111001110",
      "01011001000000101101100001001111000000000110111100010111" when "0111001111",
      "01011001001100011111011110101110111111110101011100101010" when "0111010000",
      "01011001011000010001001110011110111111100011111010101001" when "0111010001",
      "01011001100100000010110000001110111111010010010110010100" when "0111010010",
      "01011001101111110100000100011110111111000000101111101011" when "0111010011",
      "01011001111011100101001010101110111110101111000110101110" when "0111010100",
      "01011010000111010110000010111110111110011101011011011110" when "0111010101",
      "01011010010011000110101101011110111110001011101101111001" when "0111010110",
      "01011010011110110111001001111110111101111001111110000001" when "0111010111",
      "01011010101010100111011000101110111101101000001011110101" when "0111011000",
      "01011010110110010111011001001110111101010110010111010101" when "0111011001",
      "01011011000010000111001011111110111101000100100000100010" when "0111011010",
      "01011011001101110110110000011110111100110010100111011011" when "0111011011",
      "01011011011001100110000110111110111100100000101100000001" when "0111011100",
      "01011011100101010101001111011110111100001110101110010011" when "0111011101",
      "01011011110001000100001001101110111011111100101110010001" when "0111011110",
      "01011011111100110010110101111110111011101010101011111101" when "0111011111",
      "01011100001000100001010011101110111011011000100111010100" when "0111100000",
      "01011100010100001111100011101110111011000110100000011001" when "0111100001",
      "01011100011111111101100101001110111010110100010111001010" when "0111100010",
      "01011100101011101011011000011110111010100010001011101000" when "0111100011",
      "01011100110111011000111101001110111010001111111101110011" when "0111100100",
      "01011101000011000110010011111110111001111101101101101010" when "0111100101",
      "01011101001110110011011100001110111001101011011011001111" when "0111100110",
      "01011101011010100000010110001110111001011001000110100000" when "0111100111",
      "01011101100110001101000001101110111001000110101111011111" when "0111101000",
      "01011101110001111001011110101110111000110100010110001010" when "0111101001",
      "01011101111101100101101101011110111000100001111010100011" when "0111101010",
      "01011110001001010001101101011110111000001111011100101000" when "0111101011",
      "01011110010100111101011111001110110111111100111100011011" when "0111101100",
      "01011110100000101001000010001110110111101010011001111011" when "0111101101",
      "01011110101100010100010110101110110111010111110101001000" when "0111101110",
      "01011110110111111111011100011110110111000101001110000010" when "0111101111",
      "01011111000011101010010011101110110110110010100100101010" when "0111110000",
      "01011111001111010100111100011110110110011111111000111111" when "0111110001",
      "01011111011010111111010110001110110110001101001011000010" when "0111110010",
      "01011111100110101001100001011110110101111010011010110010" when "0111110011",
      "01011111110010010011011101111110110101100111101000010000" when "0111110100",
      "01011111111101111101001011101110110101010100110011011011" when "0111110101",
      "01100000001001100110101010011110110101000001111100010011" when "0111110110",
      "01100000010101001111111010011110110100101111000010111010" when "0111110111",
      "01100000100000111000111011101110110100011100000111001110" when "0111111000",
      "01100000101100100001101101111110110100001001001001010000" when "0111111001",
      "01100000111000001010010001011110110011110110001000111111" when "0111111010",
      "01100001000011110010100101111110110011100011000110011101" when "0111111011",
      "01100001001111011010101011011110110011010000000001101000" when "0111111100",
      "01100001011011000010100001111110110010111100111010100001" when "0111111101",
      "01100001100110101010001001011110110010101001110001001000" when "0111111110",
      "01100001110010010001100001101110110010010110100101011110" when "0111111111",
      "01100001111101111000101011001110110010000011010111100001" when "1000000000",
      "01100010001001011111100101001110110001110000000111010010" when "1000000001",
      "01100010010101000110010000011110110001011100110100110010" when "1000000010",
      "01100010100000101100101100011110110001001001011111111111" when "1000000011",
      "01100010101100010010111001001110110000110110001000111011" when "1000000100",
      "01100010110111111000110110101110110000100010101111100110" when "1000000101",
      "01100011000011011110100100111110110000001111010011111110" when "1000000110",
      "01100011001111000100000011111110101111111011110110000101" when "1000000111",
      "01100011011010101001010011011110101111101000010101111011" when "1000001000",
      "01100011100110001110010011111110101111010100110011011111" when "1000001001",
      "01100011110001110011000100111110101111000001001110110001" when "1000001010",
      "01100011111101010111100110011110101110101101100111110010" when "1000001011",
      "01100100001000111011111000101110101110011001111110100010" when "1000001100",
      "01100100010100011111111011011110101110000110010011000000" when "1000001101",
      "01100100100000000011101110101110101101110010100101001101" when "1000001110",
      "01100100101011100111010010101110101101011110110101001001" when "1000001111",
      "01100100110111001010100110111110101101001011000010110011" when "1000010000",
      "01100101000010101101101011011110101100110111001110001101" when "1000010001",
      "01100101001110010000100000101110101100100011010111010101" when "1000010010",
      "01100101011001110011000110001110101100001111011110001100" when "1000010011",
      "01100101100101010101011100001110101011111011100010110011" when "1000010100",
      "01100101110000110111100010001110101011100111100101001000" when "1000010101",
      "01100101111100011001011000111110101011010011100101001100" when "1000010110",
      "01100110000111111010111111101110101010111111100011000000" when "1000010111",
      "01100110010011011100010110101110101010101011011110100011" when "1000011000",
      "01100110011110111101011101111110101010010111010111110101" when "1000011001",
      "01100110101010011110010101011110101010000011001110110110" when "1000011010",
      "01100110110101111110111100111110101001101111000011100111" when "1000011011",
      "01100111000001011111010100111110101001011010110110000111" when "1000011100",
      "01100111001100111111011100101110101001000110100110010110" when "1000011101",
      "01100111011000011111010100101110101000110010010100010101" when "1000011110",
      "01100111100011111110111100101110101000011110000000000100" when "1000011111",
      "01100111101111011110010100101110101000001001101001100010" when "1000100000",
      "01100111111010111101011100111110100111110101010000110000" when "1000100001",
      "01101000000110011100010100111110100111100000110101101101" when "1000100010",
      "01101000010001111010111100111110100111001100011000011010" when "1000100011",
      "01101000011101011001010100101110100110110111111000110111" when "1000100100",
      "01101000101000110111011100101110100110100011010111000100" when "1000100101",
      "01101000110100010101010100001110100110001110110011000001" when "1000100110",
      "01101000111111110010111011101110100101111010001100101101" when "1000100111",
      "01101001001011010000010010111110100101100101100100001010" when "1000101000",
      "01101001010110101101011010001110100101010000111001010110" when "1000101001",
      "01101001100010001010010000111110100100111100001100010011" when "1000101010",
      "01101001101101100110110111011110100100100111011101000000" when "1000101011",
      "01101001111001000011001101101110100100010010101011011101" when "1000101100",
      "01101010000100011111010011101110100011111101110111101010" when "1000101101",
      "01101010001111111011001001001110100011101001000001101000" when "1000101110",
      "01101010011011010110101110011110100011010100001001010101" when "1000101111",
      "01101010100110110010000011001110100010111111001110110100" when "1000110000",
      "01101010110010001101000111101110100010101010010010000010" when "1000110001",
      "01101010111101100111111011011110100010010101010011000001" when "1000110010",
      "01101011001001000010011110101110100010000000010001110001" when "1000110011",
      "01101011010100011100110001101110100001101011001110010001" when "1000110100",
      "01101011011111110110110011111110100001010110001000100010" when "1000110101",
      "01101011101011010000100101101110100001000001000000100100" when "1000110110",
      "01101011110110101010000110101110100000101011110110010110" when "1000110111",
      "01101100000010000011010111001110100000010110101001111001" when "1000111000",
      "01101100001101011100010111001110100000000001011011001101" when "1000111001",
      "01101100011000110101000110001110011111101100001010010010" when "1000111010",
      "01101100100100001101100100101110011111010110110111000111" when "1000111011",
      "01101100101111100101110010011110011111000001100001101110" when "1000111100",
      "01101100111010111101101111001110011110101100001010000110" when "1000111101",
      "01101101000110010101011011011110011110010110110000001110" when "1000111110",
      "01101101010001101100110110101110011110000001010100001000" when "1000111111",
      "01101101011101000100000001001110011101101011110101110100" when "1001000000",
      "01101101101000011010111010101110011101010110010101010000" when "1001000001",
      "01101101110011110001100011001110011101000000110010011110" when "1001000010",
      "01101101111111000111111010111110011100101011001101011101" when "1001000011",
      "01101110001010011110000001101110011100010101100110001101" when "1001000100",
      "01101110010101110011110111011110011011111111111100101111" when "1001000101",
      "01101110100001001001011100001110011011101010010001000011" when "1001000110",
      "01101110101100011110101111111110011011010100100011001000" when "1001000111",
      "01101110110111110011110010101110011010111110110010111110" when "1001001000",
      "01101111000011001000100100001110011010101001000000100111" when "1001001001",
      "01101111001110011101000100101110011010010011001100000001" when "1001001010",
      "01101111011001110001010011111110011001111101010101001100" when "1001001011",
      "01101111100101000101010001111110011001100111011100001010" when "1001001100",
      "01101111110000011000111110111110011001010001100000111001" when "1001001101",
      "01101111111011101100011010011110011000111011100011011011" when "1001001110",
      "01110000000110111111100100111110011000100101100011101110" when "1001001111",
      "01110000010010010010011101111110011000001111100001110100" when "1001010000",
      "01110000011101100101000101101110010111111001011101101011" when "1001010001",
      "01110000101000110111011100001110010111100011010111010101" when "1001010010",
      "01110000110100001001100001001110010111001101001110110001" when "1001010011",
      "01110000111111011011010100111110010110110111000011111111" when "1001010100",
      "01110001001010101100110111001110010110100000110110111111" when "1001010101",
      "01110001010101111110000111111110010110001010100111110010" when "1001010110",
      "01110001100001001111000111001110010101110100010110010111" when "1001010111",
      "01110001101100011111110100111110010101011110000010101110" when "1001011000",
      "01110001110111110000010001001110010101000111101100111001" when "1001011001",
      "01110010000011000000011011111110010100110001010100110101" when "1001011010",
      "01110010001110010000010101001110010100011010111010100101" when "1001011011",
      "01110010011001011111111100101110010100000100011110000111" when "1001011100",
      "01110010100100101111010010011110010011101101111111011011" when "1001011101",
      "01110010101111111110010110101110010011010111011110100011" when "1001011110",
      "01110010111011001101001001001110010011000000111011011101" when "1001011111",
      "01110011000110011011101001111110010010101010010110001010" when "1001100000",
      "01110011010001101001111000111110010010010011101110101010" when "1001100001",
      "01110011011100110111110110001110010001111101000100111110" when "1001100010",
      "01110011101000000101100001101110010001100110011001000100" when "1001100011",
      "01110011110011010010111011001110010001001111101010111101" when "1001100100",
      "01110011111110100000000011001110010000111000111010101010" when "1001100101",
      "01110100001001101100111000111110010000100010001000001001" when "1001100110",
      "01110100010100111001011100111110010000001011010011011100" when "1001100111",
      "01110100100000000101101110111110001111110100011100100011" when "1001101000",
      "01110100101011010001101110111110001111011101100011011101" when "1001101001",
      "01110100110110011101011100111110001111000110101000001010" when "1001101010",
      "01110101000001101000111001001110001110101111101010101010" when "1001101011",
      "01110101001100110100000011001110001110011000101010111111" when "1001101100",
      "01110101010111111110111010111110001110000001101001000110" when "1001101101",
      "01110101100011001001100000111110001101101010100101000010" when "1001101110",
      "01110101101110010011110100011110001101010011011110110001" when "1001101111",
      "01110101111001011101110110001110001100111100010110010100" when "1001110000",
      "01110110000100100111100101011110001100100101001011101011" when "1001110001",
      "01110110001111110001000010101110001100001101111110110110" when "1001110010",
      "01110110011010111010001101011110001011110110101111110100" when "1001110011",
      "01110110100110000011000110001110001011011111011110100111" when "1001110100",
      "01110110110001001011101100011110001011001000001011001110" when "1001110101",
      "01110110111100010100000000011110001010110000110101101000" when "1001110110",
      "01110111000111011100000010001110001010011001011101110111" when "1001110111",
      "01110111010010100011110001101110001010000010000011111010" when "1001111000",
      "01110111011101101011001110011110001001101010100111110010" when "1001111001",
      "01110111101000110010011001001110001001010011001001011110" when "1001111010",
      "01110111110011111001010001001110001000111011101000111110" when "1001111011",
      "01110111111110111111110110101110001000100100000110010010" when "1001111100",
      "01111000001010000110001001111110001000001100100001011100" when "1001111101",
      "01111000010101001100001010011110000111110100111010011001" when "1001111110",
      "01111000100000010001111000011110000111011101010001001100" when "1001111111",
      "01111000101011010111010011101110000111000101100101110011" when "1010000000",
      "01111000110110011100011100101110000110101101111000001110" when "1010000001",
      "01111001000001100001010010101110000110010110001000011111" when "1010000010",
      "01111001001100100101110110001110000101111110010110100100" when "1010000011",
      "01111001010111101010000111001110000101100110100010011111" when "1010000100",
      "01111001100010101110000101001110000101001110101100001110" when "1010000101",
      "01111001101101110001110000101110000100110110110011110010" when "1010000110",
      "01111001111000110101001001001110000100011110111001001011" when "1010000111",
      "01111010000011111000001110111110000100000110111100011010" when "1010001000",
      "01111010001110111011000001111110000011101110111101011101" when "1010001001",
      "01111010011001111101100001111110000011010110111100010110" when "1010001010",
      "01111010100100111111101111001110000010111110111001000101" when "1010001011",
      "01111010110000000001101001101110000010100110110011101000" when "1010001100",
      "01111010111011000011010000111110000010001110101100000001" when "1010001101",
      "01111011000110000100100101011110000001110110100010010000" when "1010001110",
      "01111011010001000101100110111110000001011110010110010100" when "1010001111",
      "01111011011100000110010101011110000001000110001000001101" when "1010010000",
      "01111011100111000110110000111110000000101101110111111100" when "1010010001",
      "01111011110010000110111001001110000000010101100101100001" when "1010010010",
      "01111011111101000110101110011101111111111101010000111100" when "1010010011",
      "01111100001000000110010000101101111111100100111010001101" when "1010010100",
      "01111100010011000101011111101101111111001100100001010011" when "1010010101",
      "01111100011110000100011011011101111110110100000110010000" when "1010010110",
      "01111100101001000011000100001101111110011011101001000010" when "1010010111",
      "01111100110100000001011001101101111110000011001001101011" when "1010011000",
      "01111100111110111111011011111101111101101010101000001001" when "1010011001",
      "01111101001001111101001010101101111101010010000100011110" when "1010011010",
      "01111101010100111010100110011101111100111001011110101001" when "1010011011",
      "01111101011111110111101110101101111100100000110110101011" when "1010011100",
      "01111101101010110100100011011101111100001000001100100010" when "1010011101",
      "01111101110101110001000101001101111011101111100000010000" when "1010011110",
      "01111110000000101101010011001101111011010110110001110101" when "1010011111",
      "01111110001011101001001101111101111010111110000001010000" when "1010100000",
      "01111110010110100100110101001101111010100101001110100010" when "1010100001",
      "01111110100001100000001000111101111010001100011001101011" when "1010100010",
      "01111110101100011011001001001101111001110011100010101010" when "1010100011",
      "01111110110111010101110101111101111001011010101001100000" when "1010100100",
      "01111111000010010000001111001101111001000001101110001100" when "1010100101",
      "01111111001101001010010100101101111000101000110000110000" when "1010100110",
      "01111111011000000100000110101101111000001111110001001011" when "1010100111",
      "01111111100010111101100100111101110111110110101111011100" when "1010101000",
      "01111111101101110110101111101101110111011101101011100101" when "1010101001",
      "01111111111000101111100110011101110111000100100101100101" when "1010101010",
      "10000000000011101000001001101101110110101011011101011100" when "1010101011",
      "10000000001110100000011001001101110110010010010011001011" when "1010101100",
      "10000000011001011000010100111101110101111001000110110000" when "1010101101",
      "10000000100100001111111100101101110101011111111000001101" when "1010101110",
      "10000000101111000111010000111101110101000110100111100010" when "1010101111",
      "10000000111001111110010001001101110100101101010100101110" when "1010110000",
      "10000001000100110100111101011101110100010011111111110001" when "1010110001",
      "10000001001111101011010101111101110011111010101000101101" when "1010110010",
      "10000001011010100001011010011101110011100001001111011111" when "1010110011",
      "10000001100101010111001010111101110011000111110100001010" when "1010110100",
      "10000001110000001100100111011101110010101110010110101101" when "1010110101",
      "10000001111011000001101111111101110010010100110111000111" when "1010110110",
      "10000010000101110110100100011101110001111011010101011001" when "1010110111",
      "10000010010000101011000100111101110001100001110001100011" when "1010111000",
      "10000010011011011111010001011101110001001000001011100110" when "1010111001",
      "10000010100110010011001001101101110000101110100011100000" when "1010111010",
      "10000010110001000110101101101101110000010100111001010011" when "1010111011",
      "10000010111011111001111101101101101111111011001100111110" when "1010111100",
      "10000011000110101100111001011101101111100001011110100001" when "1010111101",
      "10000011010001011111100000111101101111000111101101111100" when "1010111110",
      "10000011011100010001110100001101101110101101111011010000" when "1010111111",
      "10000011100111000011110011001101101110010100000110011101" when "1011000000",
      "10000011110001110101011101111101101101111010001111100010" when "1011000001",
      "10000011111100100110110100011101101101100000010110011111" when "1011000010",
      "10000100000111010111110110011101101101000110011011010110" when "1011000011",
      "10000100010010001000100100001101101100101100011110000101" when "1011000100",
      "10000100011100111000111101011101101100010010011110101101" when "1011000101",
      "10000100100111101001000010001101101011111000011101001101" when "1011000110",
      "10000100110010011000110010101101101011011110011001100111" when "1011000111",
      "10000100111101001000001110101101101011000100010011111010" when "1011001000",
      "10000101000111110111010101111101101010101010001100000101" when "1011001001",
      "10000101010010100110001000111101101010010000000010001010" when "1011001010",
      "10000101011101010100100111001101101001110101110110001000" when "1011001011",
      "10000101101000000010110000111101101001011011100111111111" when "1011001100",
      "10000101110010110000100110001101101001000001010111110000" when "1011001101",
      "10000101111101011110000110101101101000100111000101011010" when "1011001110",
      "10000110001000001011010010101101101000001100110000111101" when "1011001111",
      "10000110010010111000001001101101100111110010011010011010" when "1011010000",
      "10000110011101100100101100001101100111011000000001110000" when "1011010001",
      "10000110101000010000111001111101100110111101100111000000" when "1011010010",
      "10000110110010111100110010111101100110100011001010001010" when "1011010011",
      "10000110111101101000010111001101100110001000101011001101" when "1011010100",
      "10000111001000010011100110011101100101101110001010001011" when "1011010101",
      "10000111010010111110100000111101100101010011100111000010" when "1011010110",
      "10000111011101101001000110101101100100111001000001110011" when "1011010111",
      "10000111101000010011010111011101100100011110011010011110" when "1011011000",
      "10000111110010111101010011011101100100000011110001000011" when "1011011001",
      "10000111111101100110111010001101100011101001000101100010" when "1011011010",
      "10001000001000010000001100001101100011001110010111111100" when "1011011011",
      "10001000010010111001001001001101100010110011101000010000" when "1011011100",
      "10001000011101100001110001001101100010011000110110011110" when "1011011101",
      "10001000101000001010000011111101100001111110000010100110" when "1011011110",
      "10001000110010110010000001111101100001100011001100101001" when "1011011111",
      "10001000111101011001101010011101100001001000010100100111" when "1011100000",
      "10001001001000000000111110001101100000101101011010011111" when "1011100001",
      "10001001010010100111111100101101100000010010011110010001" when "1011100010",
      "10001001011101001110100101111101011111110111011111111111" when "1011100011",
      "10001001100111110100111001111101011111011100011111100111" when "1011100100",
      "10001001110010011010111000111101011111000001011101001010" when "1011100101",
      "10001001111101000000100010011101011110100110011000101000" when "1011100110",
      "10001010000111100101110110111101011110001011010010000001" when "1011100111",
      "10001010010010001010110101111101011101110000001001010101" when "1011101000",
      "10001010011100101111011111101101011101010100111110100100" when "1011101001",
      "10001010100111010011110011111101011100111001110001101110" when "1011101010",
      "10001010110001110111110010111101011100011110100010110011" when "1011101011",
      "10001010111100011011011100101101011100000011010001110100" when "1011101100",
      "10001011000110111110110000101101011011100111111110110000" when "1011101101",
      "10001011010001100001101111011101011011001100101001101000" when "1011101110",
      "10001011011100000100011000101101011010110001010010011011" when "1011101111",
      "10001011100110100110101100011101011010010101111001001010" when "1011110000",
      "10001011110001001000101010101101011001111010011101110100" when "1011110001",
      "10001011111011101010010011011101011001011111000000011010" when "1011110010",
      "10001100000110001011100110011101011001000011100000111100" when "1011110011",
      "10001100010000101100100011111101011000100111111111011001" when "1011110100",
      "10001100011011001101001011101101011000001100011011110011" when "1011110101",
      "10001100100101101101011101111101010111110000110110001000" when "1011110110",
      "10001100110000001101011010011101010111010101001110011010" when "1011110111",
      "10001100111010101101000001001101010110111001100100100111" when "1011111000",
      "10001101000101001100010010001101010110011101111000110001" when "1011111001",
      "10001101001111101011001101101101010110000010001010110111" when "1011111010",
      "10001101011010001001110011001101010101100110011010111001" when "1011111011",
      "10001101100100101000000010111101010101001010101000111000" when "1011111100",
      "10001101101111000101111100101101010100101110110100110011" when "1011111101",
      "10001101111001100011100000101101010100010010111110101010" when "1011111110",
      "10001110000100000000101110111101010011110111000110011110" when "1011111111",
      "10001110001110011101100111001101010011011011001100001111" when "1100000000",
      "10001110011000111010001001011101010010111111001111111101" when "1100000001",
      "10001110100011010110010101111101010010100011010001100111" when "1100000010",
      "10001110101101110010001100001101010010000111010001001110" when "1100000011",
      "10001110111000001101101100101101010001101011001110110010" when "1100000100",
      "10001111000010101000110110111101010001001111001010010011" when "1100000101",
      "10001111001101000011101011001101010000110011000011110001" when "1100000110",
      "10001111010111011110001001011101010000010110111011001100" when "1100000111",
      "10001111100001111000010001011101001111111010110000100100" when "1100001000",
      "10001111101100010010000011011101001111011110100011111010" when "1100001001",
      "10001111110110101011011111001101001111000010010101001100" when "1100001010",
      "10010000000001000100100100101101001110100110000100011100" when "1100001011",
      "10010000001011011101010100001101001110001001110001101010" when "1100001100",
      "10010000010101110101101101001101001101101101011100110101" when "1100001101",
      "10010000100000001101110000001101001101010001000101111110" when "1100001110",
      "10010000101010100101011100101101001100110100101101000100" when "1100001111",
      "10010000110100111100110011001101001100011000010010001000" when "1100010000",
      "10010000111111010011110010111101001011111011110101001010" when "1100010001",
      "10010001001001101010011100101101001011011111010110001010" when "1100010010",
      "10010001010100000000101111111101001011000010110101000111" when "1100010011",
      "10010001011110010110101100101101001010100110010010000011" when "1100010100",
      "10010001101000101100010011001101001010001001101100111101" when "1100010101",
      "10010001110011000001100010111101001001101101000101110101" when "1100010110",
      "10010001111101010110011100011101001001010000011100101011" when "1100010111",
      "10010010000111101010111111011101001000110011110001011111" when "1100011000",
      "10010010010001111111001011101101001000010111000100010010" when "1100011001",
      "10010010011100010011000001101101000111111010010101000011" when "1100011010",
      "10010010100110100110100000111101000111011101100011110010" when "1100011011",
      "10010010110000111001101001011101000111000000110000100000" when "1100011100",
      "10010010111011001100011011011101000110100011111011001101" when "1100011101",
      "10010011000101011110110110111101000110000111000011111000" when "1100011110",
      "10010011001111110000111011011101000101101010001010100010" when "1100011111",
      "10010011011010000010101001011101000101001101001111001011" when "1100100000",
      "10010011100100010100000000101101000100110000010001110011" when "1100100001",
      "10010011101110100101000001001101000100010011010010011010" when "1100100010",
      "10010011111000110101101010111101000011110110010000111111" when "1100100011",
      "10010100000011000101111101101101000011011001001101100100" when "1100100100",
      "10010100001101010101111001111101000010111100001000001000" when "1100100101",
      "10010100010111100101011110111101000010011111000000101100" when "1100100110",
      "10010100100001110100101101011101000010000001110111001110" when "1100100111",
      "10010100101100000011100100101101000001100100101011110000" when "1100101000",
      "10010100110110010010000101001101000001000111011110010010" when "1100101001",
      "10010101000000100000001110101101000000101010001110110011" when "1100101010",
      "10010101001010101110000001011101000000001100111101010011" when "1100101011",
      "10010101010100111011011100111100111111101111101001110100" when "1100101100",
      "10010101011111001000100001011100111111010010010100010100" when "1100101101",
      "10010101101001010101001110111100111110110100111100110011" when "1100101110",
      "10010101110011100001100101001100111110010111100011010011" when "1100101111",
      "10010101111101101101100100101100111101111010000111110011" when "1100110000",
      "10010110000111111001001100101100111101011100101010010010" when "1100110001",
      "10010110010010000100011101101100111100111111001010110010" when "1100110010",
      "10010110011100001111010111101100111100100001101001010010" when "1100110011",
      "10010110100110011001111010001100111100000100000101110010" when "1100110100",
      "10010110110000100100000101101100111011100110100000010010" when "1100110101",
      "10010110111010101101111001111100111011001000111000110011" when "1100110110",
      "10010111000100110111010110101100111010101011001111010100" when "1100110111",
      "10010111001111000000011100011100111010001101100011110110" when "1100111000",
      "10010111011001001001001010101100111001101111110110011000" when "1100111001",
      "10010111100011010001100001011100111001010010000110111011" when "1100111010",
      "10010111101101011001100001001100111000110100010101011111" when "1100111011",
      "10010111110111100001001001001100111000010110100010000100" when "1100111100",
      "10011000000001101000011001111100110111111000101100101001" when "1100111101",
      "10011000001011101111010011001100110111011010110101001111" when "1100111110",
      "10011000010101110101110101001100110110111100111011110111" when "1100111111",
      "10011000011111111011111111011100110110011111000000011111" when "1101000000",
      "10011000101010000001110010001100110110000001000011001001" when "1101000001",
      "10011000110100000111001101011100110101100011000011110100" when "1101000010",
      "10011000111110001100010001001100110101000101000010100000" when "1101000011",
      "10011001001000010000111101011100110100100110111111001101" when "1101000100",
      "10011001010010010101010001111100110100001000111001111100" when "1101000101",
      "10011001011100011001001110101100110011101010110010101101" when "1101000110",
      "10011001100110011100110011111100110011001100101001011111" when "1101000111",
      "10011001110000100000000001011100110010101110011110010011" when "1101001000",
      "10011001111010100010110111001100110010010000010001001000" when "1101001001",
      "10011010000100100101010101001100110001110010000001111111" when "1101001010",
      "10011010001110100111011011101100110001010011110000111001" when "1101001011",
      "10011010011000101001001010001100110000110101011101110100" when "1101001100",
      "10011010100010101010100000111100110000010111001000110001" when "1101001101",
      "10011010101100101011011111101100101111111000110001110000" when "1101001110",
      "10011010110110101100000110101100101111011010011000110010" when "1101001111",
      "10011011000000101100010101111100101110111011111101110110" when "1101010000",
      "10011011001010101100001101001100101110011101100000111100" when "1101010001",
      "10011011010100101011101100011100101101111111000010000100" when "1101010010",
      "10011011011110101010110011101100101101100000100001001111" when "1101010011",
      "10011011101000101001100011001100101101000001111110011101" when "1101010100",
      "10011011110010100111111010101100101100100011011001101101" when "1101010101",
      "10011011111100100101111001111100101100000100110011000000" when "1101010110",
      "10011100000110100011100001001100101011100110001010010101" when "1101010111",
      "10011100010000100000110000011100101011000111011111101110" when "1101011000",
      "10011100011010011101100111101100101010101000110011001001" when "1101011001",
      "10011100100100011010000110101100101010001010000100100111" when "1101011010",
      "10011100101110010110001101011100101001101011010100001001" when "1101011011",
      "10011100111000010001111100001100101001001100100001101101" when "1101011100",
      "10011101000010001101010010101100101000101101101101010101" when "1101011101",
      "10011101001100001000010000111100101000001110110111000000" when "1101011110",
      "10011101010110000010110111001100100111101111111110101110" when "1101011111",
      "10011101011111111101000100111100100111010001000100100000" when "1101100000",
      "10011101101001110110111010011100100110110010001000010110" when "1101100001",
      "10011101110011110000010111011100100110010011001010001110" when "1101100010",
      "10011101111101101001011100011100100101110100001010001011" when "1101100011",
      "10011110000111100010001000111100100101010101001000001011" when "1101100100",
      "10011110010001011010011100111100100100110110000100001111" when "1101100101",
      "10011110011011010010011000101100100100010110111110010111" when "1101100110",
      "10011110100101001001111011111100100011110111110110100011" when "1101100111",
      "10011110101111000001000110101100100011011000101100110011" when "1101101000",
      "10011110111000110111111001001100100010111001100001000111" when "1101101001",
      "10011111000010101110010010111100100010011010010011100000" when "1101101010",
      "10011111001100100100010100001100100001111011000011111100" when "1101101011",
      "10011111010110011001111100111100100001011011110010011101" when "1101101100",
      "10011111100000001111001101001100100000111100011111000010" when "1101101101",
      "10011111101010000100000100101100100000011101001001101100" when "1101101110",
      "10011111110011111000100011101100011111111101110010011011" when "1101101111",
      "10011111111101101100101010001100011111011110011001001101" when "1101110000",
      "10100000000111100000010111101100011110111110111110000101" when "1101110001",
      "10100000010001010011101100101100011110011111100001000010" when "1101110010",
      "10100000011011000110101000111100011110000000000010000011" when "1101110011",
      "10100000100100111001001100011100011101100000100001001001" when "1101110100",
      "10100000101110101011010111001100011101000000111110010100" when "1101110101",
      "10100000111000011101001001001100011100100001011001100101" when "1101110110",
      "10100001000010001110100010001100011100000001110010111010" when "1101110111",
      "10100001001011111111100010101100011011100010001010010101" when "1101111000",
      "10100001010101110000001010001100011011000010011111110101" when "1101111001",
      "10100001011111100000011000101100011010100010110011011011" when "1101111010",
      "10100001101001010000001110011100011010000011000101000110" when "1101111011",
      "10100001110010111111101010111100011001100011010100110110" when "1101111100",
      "10100001111100101110101110111100011001000011100010101100" when "1101111101",
      "10100010000110011101011001101100011000100011101110101000" when "1101111110",
      "10100010010000001011101011011100011000000011111000101010" when "1101111111",
      "10100010011001111001100100001100010111100100000000110001" when "1110000000",
      "10100010100011100111000011111100010111000100000110111111" when "1110000001",
      "10100010101101010100001010101100010110100100001011010010" when "1110000010",
      "10100010110111000000111000001100010110000100001101101011" when "1110000011",
      "10100011000000101101001100101100010101100100001110001011" when "1110000100",
      "10100011001010011001001000001100010101000100001100110001" when "1110000101",
      "10100011010100000100101010001100010100100100001001011101" when "1110000110",
      "10100011011101101111110011001100010100000100000100010000" when "1110000111",
      "10100011100111011010100011001100010011100011111101001001" when "1110001000",
      "10100011110001000100111001101100010011000011110100001000" when "1110001001",
      "10100011111010101110110110111100010010100011101001001111" when "1110001010",
      "10100100000100011000011010111100010010000011011100011100" when "1110001011",
      "10100100001110000001100101101100010001100011001101101111" when "1110001100",
      "10100100010111101010010110111100010001000010111101001010" when "1110001101",
      "10100100100001010010101111001100010000100010101010101011" when "1110001110",
      "10100100101010111010101101101100010000000010010110010100" when "1110001111",
      "10100100110100100010010011001100001111100010000000000100" when "1110010000",
      "10100100111110001001011110111100001111000001100111111010" when "1110010001",
      "10100101000111110000010001011100001110100001001101111000" when "1110010010",
      "10100101010001010110101010001100001110000000110001111110" when "1110010011",
      "10100101011010111100101001101100001101100000010100001011" when "1110010100",
      "10100101100100100010001111101100001100111111110100011111" when "1110010101",
      "10100101101110000111011100001100001100011111010010111011" when "1110010110",
      "10100101110111101100001110111100001011111110101111011110" when "1110010111",
      "10100110000001010000101000011100001011011110001010001001" when "1110011000",
      "10100110001010110100100111111100001010111101100010111100" when "1110011001",
      "10100110010100011000001110001100001010011100111001110111" when "1110011010",
      "10100110011101111011011010011100001001111100001110111010" when "1110011011",
      "10100110100111011110001101001100001001011011100010000101" when "1110011100",
      "10100110110001000000100110001100001000111010110011011000" when "1110011101",
      "10100110111010100010100101101100001000011010000010110011" when "1110011110",
      "10100111000100000100001011001100000111111001010000010110" when "1110011111",
      "10100111001101100101010110111100000111011000011100000010" when "1110100000",
      "10100111010111000110001001001100000110110111100101110110" when "1110100001",
      "10100111100000100110100001011100000110010110101101110011" when "1110100010",
      "10100111101010000110011111101100000101110101110011111000" when "1110100011",
      "10100111110011100110000100001100000101010100111000000110" when "1110100100",
      "10100111111101000101001110111100000100110011111010011101" when "1110100101",
      "10101000000110100011111111101100000100010010111010111100" when "1110100110",
      "10101000010000000010010110101100000011110001111001100100" when "1110100111",
      "10101000011001100000010011011100000011010000110110010110" when "1110101000",
      "10101000100010111101110110011100000010101111110001010000" when "1110101001",
      "10101000101100011010111111011100000010001110101010010100" when "1110101010",
      "10101000110101110111101110001100000001101101100001100001" when "1110101011",
      "10101000111111010100000011001100000001001100010110110111" when "1110101100",
      "10101001001000101111111101111100000000101011001010010110" when "1110101101",
      "10101001010010001011011110101100000000001001111011111111" when "1110101110",
      "10101001011011100110100101011011111111101000101011110010" when "1110101111",
      "10101001100101000001010001111011111111000111011001101110" when "1110110000",
      "10101001101110011011100100001011111110100110000101110011" when "1110110001",
      "10101001110111110101011100011011111110000100110000000011" when "1110110010",
      "10101010000001001110111010011011111101100011011000011101" when "1110110011",
      "10101010001010100111111110001011111101000001111111000000" when "1110110100",
      "10101010010100000000100111101011111100100000100011101101" when "1110110101",
      "10101010011101011000110110111011111011111111000110100101" when "1110110110",
      "10101010100110110000101011111011111011011101100111100111" when "1110110111",
      "10101010110000001000000110101011111010111100000110110010" when "1110111000",
      "10101010111001011111000110111011111010011010100100001001" when "1110111001",
      "10101011000010110101101100111011111001111000111111101001" when "1110111010",
      "10101011001100001011111000011011111001010111011001010101" when "1110111011",
      "10101011010101100001101001101011111000110101110001001011" when "1110111100",
      "10101011011110110111000000011011111000010100000111001011" when "1110111101",
      "10101011101000001011111100111011110111110010011011010110" when "1110111110",
      "10101011110001100000011110101011110111010000101101101100" when "1110111111",
      "10101011111010110100100110001011110110101110111110001101" when "1111000000",
      "10101100000100001000010010111011110110001101001100111001" when "1111000001",
      "10101100001101011011100101001011110101101011011001110000" when "1111000010",
      "10101100010110101110011100111011110101001001100100110011" when "1111000011",
      "10101100100000000000111010001011110100100111101110000000" when "1111000100",
      "10101100101001010010111100111011110100000101110101011001" when "1111000101",
      "10101100110010100100100100101011110011100011111010111101" when "1111000110",
      "10101100111011110101110010001011110011000001111110101101" when "1111000111",
      "10101101000101000110100100101011110010100000000000101000" when "1111001000",
      "10101101001110010110111100101011110001111110000000101111" when "1111001001",
      "10101101010111100110111001111011110001011011111111000001" when "1111001010",
      "10101101100000110110011100011011110000111001111011100000" when "1111001011",
      "10101101101010000101100100001011110000010111110110001010" when "1111001100",
      "10101101110011010100010001001011101111110101101111000000" when "1111001101",
      "10101101111100100010100011011011101111010011100110000011" when "1111001110",
      "10101110000101110000011010101011101110110001011011010001" when "1111001111",
      "10101110001110111101110111001011101110001111001110101100" when "1111010000",
      "10101110011000001010111000111011101101101101000000010011" when "1111010001",
      "10101110100001010111011111101011101101001010110000000110" when "1111010010",
      "10101110101010100011101011011011101100101000011110000110" when "1111010011",
      "10101110110011101111011100011011101100000110001010010010" when "1111010100",
      "10101110111100111010110010001011101011100011110100101011" when "1111010101",
      "10101111000110000101101101001011101011000001011101010001" when "1111010110",
      "10101111001111010000001101001011101010011111000100000100" when "1111010111",
      "10101111011000011010010010001011101001111100101001000011" when "1111011000",
      "10101111100001100011111011111011101001011010001100010000" when "1111011001",
      "10101111101010101101001010111011101000110111101101101001" when "1111011010",
      "10101111110011110101111110011011101000010101001101010000" when "1111011011",
      "10101111111100111110010111001011100111110010101011000011" when "1111011100",
      "10110000000110000110010100101011100111010000000111000100" when "1111011101",
      "10110000001111001101110110111011100110101101100001010011" when "1111011110",
      "10110000011000010100111110001011100110001010111001101111" when "1111011111",
      "10110000100001011011101010001011100101101000010000011000" when "1111100000",
      "10110000101010100001111010101011100101000101100101001111" when "1111100001",
      "10110000110011100111110000001011100100100010111000010100" when "1111100010",
      "10110000111100101101001010011011100100000000001001100111" when "1111100011",
      "10110001000101110010001001011011100011011101011001000111" when "1111100100",
      "10110001001110110110101100111011100010111010100110110110" when "1111100101",
      "10110001010111111010110101001011100010010111110010110010" when "1111100110",
      "10110001100000111110100010001011100001110100111100111101" when "1111100111",
      "10110001101010000001110011101011100001010010000101010110" when "1111101000",
      "10110001110011000100101001111011100000101111001011111101" when "1111101001",
      "10110001111100000111000100101011100000001100010000110011" when "1111101010",
      "10110010000101001001000011111011011111101001010011110111" when "1111101011",
      "10110010001110001010100111111011011111000110010101001001" when "1111101100",
      "10110010010111001011110000001011011110100011010100101011" when "1111101101",
      "10110010100000001100011100111011011110000000010010011011" when "1111101110",
      "10110010101001001100101110011011011101011101001110011001" when "1111101111",
      "10110010110010001100100100001011011100111010001000100111" when "1111110000",
      "10110010111011001011111110011011011100010111000001000100" when "1111110001",
      "10110011000100001010111100111011011011110011110111101111" when "1111110010",
      "10110011001101001001011111111011011011010000101100101010" when "1111110011",
      "10110011010110000111100111001011011010101101011111110100" when "1111110100",
      "10110011011111000101010010111011011010001010010001001110" when "1111110101",
      "10110011101000000010100010111011011001100111000000110110" when "1111110110",
      "10110011110000111111010111011011011001000011101110101111" when "1111110111",
      "10110011111001111011101111111011011000100000011010110110" when "1111111000",
      "10110100000010110111101100101011010111111101000101001110" when "1111111001",
      "10110100001011110011001101111011010111011001101101110101" when "1111111010",
      "10110100010100101110010011001011010110110110010100101100" when "1111111011",
      "10110100011101101000111100101011010110010010111001110011" when "1111111100",
      "10110100100110100011001010011011010101101111011101001010" when "1111111101",
      "10110100101111011100111100001011010101001011111110110001" when "1111111110",
      "10110100111000010110010010001011010100101000011110101000" when "1111111111",
      "--------------------------------------------------------" when others;
   Y1 <= Y0_d1; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_19_Freq200_uid39
-- VHDL generated for DummyFPGA @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X Y Cin
-- Output signals: R
--  approx. input signal timings: X: (c0, 1.700000ns)Y: (c0, 1.700000ns)Cin: (c0, 0.000000ns)
--  approx. output signal timings: R: (c0, 2.880000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_19_Freq200_uid39 is
    port (clk, rst : in std_logic;
          X : in  std_logic_vector(18 downto 0);
          Y : in  std_logic_vector(18 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(18 downto 0)   );
end entity;

architecture arch of IntAdder_19_Freq200_uid39 is
signal Rtmp :  std_logic_vector(18 downto 0);
   -- timing of Rtmp: (c0, 2.880000ns)
begin
   Rtmp <= X + Y + Cin;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          FixRealKCM_Freq200_uid6
-- VHDL generated for DummyFPGA @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: R
--  approx. input signal timings: X: (c0, 0.550000ns)
--  approx. output signal timings: R: (c0, 2.880000ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixRealKCM_Freq200_uid6 is
    port (clk, rst : in std_logic;
          X : in  std_logic_vector(15 downto 0);
          R : out  std_logic_vector(17 downto 0)   );
end entity;

architecture arch of FixRealKCM_Freq200_uid6 is
   component FixRealKCM_Freq200_uid6_T0_Freq200_uid9 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(19 downto 0)   );
   end component;

   component FixRealKCM_Freq200_uid6_T1_Freq200_uid12 is
      port ( X : in  std_logic_vector(4 downto 0);
             Y : out  std_logic_vector(14 downto 0)   );
   end component;

   component FixRealKCM_Freq200_uid6_T2_Freq200_uid15 is
      port ( X : in  std_logic_vector(5 downto 0);
             Y : out  std_logic_vector(9 downto 0)   );
   end component;

   component Compressor_23_3_Freq200_uid19 is
      port ( X1 : in  std_logic_vector(1 downto 0);
             X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_14_3_Freq200_uid35 is
      port ( X1 : in  std_logic_vector(0 downto 0);
             X0 : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component IntAdder_19_Freq200_uid39 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(18 downto 0);
             Y : in  std_logic_vector(18 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(18 downto 0)   );
   end component;

signal FixRealKCM_Freq200_uid6_A0 :  std_logic_vector(4 downto 0);
   -- timing of FixRealKCM_Freq200_uid6_A0: (c0, 0.550000ns)
signal FixRealKCM_Freq200_uid6_T0 :  std_logic_vector(19 downto 0);
   -- timing of FixRealKCM_Freq200_uid6_T0: (c0, 1.100000ns)
signal FixRealKCM_Freq200_uid6_T0_copy10 :  std_logic_vector(19 downto 0);
   -- timing of FixRealKCM_Freq200_uid6_T0_copy10: (c0, 0.550000ns)
signal bh7_w0_0 :  std_logic;
   -- timing of bh7_w0_0: (c0, 1.100000ns)
signal bh7_w1_0 :  std_logic;
   -- timing of bh7_w1_0: (c0, 1.100000ns)
signal bh7_w2_0 :  std_logic;
   -- timing of bh7_w2_0: (c0, 1.100000ns)
signal bh7_w3_0 :  std_logic;
   -- timing of bh7_w3_0: (c0, 1.100000ns)
signal bh7_w4_0 :  std_logic;
   -- timing of bh7_w4_0: (c0, 1.100000ns)
signal bh7_w5_0 :  std_logic;
   -- timing of bh7_w5_0: (c0, 1.100000ns)
signal bh7_w6_0 :  std_logic;
   -- timing of bh7_w6_0: (c0, 1.100000ns)
signal bh7_w7_0 :  std_logic;
   -- timing of bh7_w7_0: (c0, 1.100000ns)
signal bh7_w8_0 :  std_logic;
   -- timing of bh7_w8_0: (c0, 1.100000ns)
signal bh7_w9_0 :  std_logic;
   -- timing of bh7_w9_0: (c0, 1.100000ns)
signal bh7_w10_0 :  std_logic;
   -- timing of bh7_w10_0: (c0, 1.100000ns)
signal bh7_w11_0 :  std_logic;
   -- timing of bh7_w11_0: (c0, 1.100000ns)
signal bh7_w12_0 :  std_logic;
   -- timing of bh7_w12_0: (c0, 1.100000ns)
signal bh7_w13_0 :  std_logic;
   -- timing of bh7_w13_0: (c0, 1.100000ns)
signal bh7_w14_0 :  std_logic;
   -- timing of bh7_w14_0: (c0, 1.100000ns)
signal bh7_w15_0 :  std_logic;
   -- timing of bh7_w15_0: (c0, 1.100000ns)
signal bh7_w16_0 :  std_logic;
   -- timing of bh7_w16_0: (c0, 1.100000ns)
signal bh7_w17_0 :  std_logic;
   -- timing of bh7_w17_0: (c0, 1.100000ns)
signal bh7_w18_0 :  std_logic;
   -- timing of bh7_w18_0: (c0, 1.100000ns)
signal bh7_w19_0 :  std_logic;
   -- timing of bh7_w19_0: (c0, 1.100000ns)
signal FixRealKCM_Freq200_uid6_A1 :  std_logic_vector(4 downto 0);
   -- timing of FixRealKCM_Freq200_uid6_A1: (c0, 0.550000ns)
signal FixRealKCM_Freq200_uid6_T1 :  std_logic_vector(14 downto 0);
   -- timing of FixRealKCM_Freq200_uid6_T1: (c0, 1.100000ns)
signal FixRealKCM_Freq200_uid6_T1_copy13 :  std_logic_vector(14 downto 0);
   -- timing of FixRealKCM_Freq200_uid6_T1_copy13: (c0, 0.550000ns)
signal bh7_w0_1 :  std_logic;
   -- timing of bh7_w0_1: (c0, 1.100000ns)
signal bh7_w1_1 :  std_logic;
   -- timing of bh7_w1_1: (c0, 1.100000ns)
signal bh7_w2_1 :  std_logic;
   -- timing of bh7_w2_1: (c0, 1.100000ns)
signal bh7_w3_1 :  std_logic;
   -- timing of bh7_w3_1: (c0, 1.100000ns)
signal bh7_w4_1 :  std_logic;
   -- timing of bh7_w4_1: (c0, 1.100000ns)
signal bh7_w5_1 :  std_logic;
   -- timing of bh7_w5_1: (c0, 1.100000ns)
signal bh7_w6_1 :  std_logic;
   -- timing of bh7_w6_1: (c0, 1.100000ns)
signal bh7_w7_1 :  std_logic;
   -- timing of bh7_w7_1: (c0, 1.100000ns)
signal bh7_w8_1 :  std_logic;
   -- timing of bh7_w8_1: (c0, 1.100000ns)
signal bh7_w9_1 :  std_logic;
   -- timing of bh7_w9_1: (c0, 1.100000ns)
signal bh7_w10_1 :  std_logic;
   -- timing of bh7_w10_1: (c0, 1.100000ns)
signal bh7_w11_1 :  std_logic;
   -- timing of bh7_w11_1: (c0, 1.100000ns)
signal bh7_w12_1 :  std_logic;
   -- timing of bh7_w12_1: (c0, 1.100000ns)
signal bh7_w13_1 :  std_logic;
   -- timing of bh7_w13_1: (c0, 1.100000ns)
signal bh7_w14_1 :  std_logic;
   -- timing of bh7_w14_1: (c0, 1.100000ns)
signal FixRealKCM_Freq200_uid6_A2 :  std_logic_vector(5 downto 0);
   -- timing of FixRealKCM_Freq200_uid6_A2: (c0, 0.550000ns)
signal FixRealKCM_Freq200_uid6_T2 :  std_logic_vector(9 downto 0);
   -- timing of FixRealKCM_Freq200_uid6_T2: (c0, 1.150000ns)
signal FixRealKCM_Freq200_uid6_T2_copy16 :  std_logic_vector(9 downto 0);
   -- timing of FixRealKCM_Freq200_uid6_T2_copy16: (c0, 0.550000ns)
signal bh7_w0_2 :  std_logic;
   -- timing of bh7_w0_2: (c0, 1.150000ns)
signal bh7_w1_2 :  std_logic;
   -- timing of bh7_w1_2: (c0, 1.150000ns)
signal bh7_w2_2 :  std_logic;
   -- timing of bh7_w2_2: (c0, 1.150000ns)
signal bh7_w3_2 :  std_logic;
   -- timing of bh7_w3_2: (c0, 1.150000ns)
signal bh7_w4_2 :  std_logic;
   -- timing of bh7_w4_2: (c0, 1.150000ns)
signal bh7_w5_2 :  std_logic;
   -- timing of bh7_w5_2: (c0, 1.150000ns)
signal bh7_w6_2 :  std_logic;
   -- timing of bh7_w6_2: (c0, 1.150000ns)
signal bh7_w7_2 :  std_logic;
   -- timing of bh7_w7_2: (c0, 1.150000ns)
signal bh7_w8_2 :  std_logic;
   -- timing of bh7_w8_2: (c0, 1.150000ns)
signal bh7_w9_2 :  std_logic;
   -- timing of bh7_w9_2: (c0, 1.150000ns)
signal Compressor_23_3_Freq200_uid19_bh7_uid20_In0 :  std_logic_vector(2 downto 0);
   -- timing of Compressor_23_3_Freq200_uid19_bh7_uid20_In0: (c0, 1.150000ns)
signal Compressor_23_3_Freq200_uid19_bh7_uid20_In1 :  std_logic_vector(1 downto 0);
   -- timing of Compressor_23_3_Freq200_uid19_bh7_uid20_In1: (c0, 1.100000ns)
signal Compressor_23_3_Freq200_uid19_bh7_uid20_Out0 :  std_logic_vector(2 downto 0);
   -- timing of Compressor_23_3_Freq200_uid19_bh7_uid20_Out0: (c0, 1.700000ns)
signal bh7_w0_3 :  std_logic;
   -- timing of bh7_w0_3: (c0, 1.700000ns)
signal bh7_w1_3 :  std_logic;
   -- timing of bh7_w1_3: (c0, 1.700000ns)
signal bh7_w2_3 :  std_logic;
   -- timing of bh7_w2_3: (c0, 1.700000ns)
signal Compressor_23_3_Freq200_uid19_bh7_uid20_Out0_copy21 :  std_logic_vector(2 downto 0);
   -- timing of Compressor_23_3_Freq200_uid19_bh7_uid20_Out0_copy21: (c0, 1.150000ns)
signal Compressor_23_3_Freq200_uid19_bh7_uid22_In0 :  std_logic_vector(2 downto 0);
   -- timing of Compressor_23_3_Freq200_uid19_bh7_uid22_In0: (c0, 1.150000ns)
signal Compressor_23_3_Freq200_uid19_bh7_uid22_In1 :  std_logic_vector(1 downto 0);
   -- timing of Compressor_23_3_Freq200_uid19_bh7_uid22_In1: (c0, 1.100000ns)
signal Compressor_23_3_Freq200_uid19_bh7_uid22_Out0 :  std_logic_vector(2 downto 0);
   -- timing of Compressor_23_3_Freq200_uid19_bh7_uid22_Out0: (c0, 1.700000ns)
signal bh7_w2_4 :  std_logic;
   -- timing of bh7_w2_4: (c0, 1.700000ns)
signal bh7_w3_3 :  std_logic;
   -- timing of bh7_w3_3: (c0, 1.700000ns)
signal bh7_w4_3 :  std_logic;
   -- timing of bh7_w4_3: (c0, 1.700000ns)
signal Compressor_23_3_Freq200_uid19_bh7_uid22_Out0_copy23 :  std_logic_vector(2 downto 0);
   -- timing of Compressor_23_3_Freq200_uid19_bh7_uid22_Out0_copy23: (c0, 1.150000ns)
signal Compressor_23_3_Freq200_uid19_bh7_uid24_In0 :  std_logic_vector(2 downto 0);
   -- timing of Compressor_23_3_Freq200_uid19_bh7_uid24_In0: (c0, 1.150000ns)
signal Compressor_23_3_Freq200_uid19_bh7_uid24_In1 :  std_logic_vector(1 downto 0);
   -- timing of Compressor_23_3_Freq200_uid19_bh7_uid24_In1: (c0, 1.100000ns)
signal Compressor_23_3_Freq200_uid19_bh7_uid24_Out0 :  std_logic_vector(2 downto 0);
   -- timing of Compressor_23_3_Freq200_uid19_bh7_uid24_Out0: (c0, 1.700000ns)
signal bh7_w4_4 :  std_logic;
   -- timing of bh7_w4_4: (c0, 1.700000ns)
signal bh7_w5_3 :  std_logic;
   -- timing of bh7_w5_3: (c0, 1.700000ns)
signal bh7_w6_3 :  std_logic;
   -- timing of bh7_w6_3: (c0, 1.700000ns)
signal Compressor_23_3_Freq200_uid19_bh7_uid24_Out0_copy25 :  std_logic_vector(2 downto 0);
   -- timing of Compressor_23_3_Freq200_uid19_bh7_uid24_Out0_copy25: (c0, 1.150000ns)
signal Compressor_23_3_Freq200_uid19_bh7_uid26_In0 :  std_logic_vector(2 downto 0);
   -- timing of Compressor_23_3_Freq200_uid19_bh7_uid26_In0: (c0, 1.150000ns)
signal Compressor_23_3_Freq200_uid19_bh7_uid26_In1 :  std_logic_vector(1 downto 0);
   -- timing of Compressor_23_3_Freq200_uid19_bh7_uid26_In1: (c0, 1.100000ns)
signal Compressor_23_3_Freq200_uid19_bh7_uid26_Out0 :  std_logic_vector(2 downto 0);
   -- timing of Compressor_23_3_Freq200_uid19_bh7_uid26_Out0: (c0, 1.700000ns)
signal bh7_w6_4 :  std_logic;
   -- timing of bh7_w6_4: (c0, 1.700000ns)
signal bh7_w7_3 :  std_logic;
   -- timing of bh7_w7_3: (c0, 1.700000ns)
signal bh7_w8_3 :  std_logic;
   -- timing of bh7_w8_3: (c0, 1.700000ns)
signal Compressor_23_3_Freq200_uid19_bh7_uid26_Out0_copy27 :  std_logic_vector(2 downto 0);
   -- timing of Compressor_23_3_Freq200_uid19_bh7_uid26_Out0_copy27: (c0, 1.150000ns)
signal Compressor_23_3_Freq200_uid19_bh7_uid28_In0 :  std_logic_vector(2 downto 0);
   -- timing of Compressor_23_3_Freq200_uid19_bh7_uid28_In0: (c0, 1.150000ns)
signal Compressor_23_3_Freq200_uid19_bh7_uid28_In1 :  std_logic_vector(1 downto 0);
   -- timing of Compressor_23_3_Freq200_uid19_bh7_uid28_In1: (c0, 1.100000ns)
signal Compressor_23_3_Freq200_uid19_bh7_uid28_Out0 :  std_logic_vector(2 downto 0);
   -- timing of Compressor_23_3_Freq200_uid19_bh7_uid28_Out0: (c0, 1.700000ns)
signal bh7_w8_4 :  std_logic;
   -- timing of bh7_w8_4: (c0, 1.700000ns)
signal bh7_w9_3 :  std_logic;
   -- timing of bh7_w9_3: (c0, 1.700000ns)
signal bh7_w10_2 :  std_logic;
   -- timing of bh7_w10_2: (c0, 1.700000ns)
signal Compressor_23_3_Freq200_uid19_bh7_uid28_Out0_copy29 :  std_logic_vector(2 downto 0);
   -- timing of Compressor_23_3_Freq200_uid19_bh7_uid28_Out0_copy29: (c0, 1.150000ns)
signal Compressor_23_3_Freq200_uid19_bh7_uid30_In0 :  std_logic_vector(2 downto 0);
   -- timing of Compressor_23_3_Freq200_uid19_bh7_uid30_In0: (c0, 1.100000ns)
signal Compressor_23_3_Freq200_uid19_bh7_uid30_In1 :  std_logic_vector(1 downto 0);
   -- timing of Compressor_23_3_Freq200_uid19_bh7_uid30_In1: (c0, 1.100000ns)
signal Compressor_23_3_Freq200_uid19_bh7_uid30_Out0 :  std_logic_vector(2 downto 0);
   -- timing of Compressor_23_3_Freq200_uid19_bh7_uid30_Out0: (c0, 1.650000ns)
signal bh7_w10_3 :  std_logic;
   -- timing of bh7_w10_3: (c0, 1.650000ns)
signal bh7_w11_2 :  std_logic;
   -- timing of bh7_w11_2: (c0, 1.650000ns)
signal bh7_w12_2 :  std_logic;
   -- timing of bh7_w12_2: (c0, 1.650000ns)
signal Compressor_23_3_Freq200_uid19_bh7_uid30_Out0_copy31 :  std_logic_vector(2 downto 0);
   -- timing of Compressor_23_3_Freq200_uid19_bh7_uid30_Out0_copy31: (c0, 1.100000ns)
signal Compressor_23_3_Freq200_uid19_bh7_uid32_In0 :  std_logic_vector(2 downto 0);
   -- timing of Compressor_23_3_Freq200_uid19_bh7_uid32_In0: (c0, 1.100000ns)
signal Compressor_23_3_Freq200_uid19_bh7_uid32_In1 :  std_logic_vector(1 downto 0);
   -- timing of Compressor_23_3_Freq200_uid19_bh7_uid32_In1: (c0, 1.100000ns)
signal Compressor_23_3_Freq200_uid19_bh7_uid32_Out0 :  std_logic_vector(2 downto 0);
   -- timing of Compressor_23_3_Freq200_uid19_bh7_uid32_Out0: (c0, 1.650000ns)
signal bh7_w12_3 :  std_logic;
   -- timing of bh7_w12_3: (c0, 1.650000ns)
signal bh7_w13_2 :  std_logic;
   -- timing of bh7_w13_2: (c0, 1.650000ns)
signal bh7_w14_2 :  std_logic;
   -- timing of bh7_w14_2: (c0, 1.650000ns)
signal Compressor_23_3_Freq200_uid19_bh7_uid32_Out0_copy33 :  std_logic_vector(2 downto 0);
   -- timing of Compressor_23_3_Freq200_uid19_bh7_uid32_Out0_copy33: (c0, 1.100000ns)
signal Compressor_14_3_Freq200_uid35_bh7_uid36_In0 :  std_logic_vector(3 downto 0);
   -- timing of Compressor_14_3_Freq200_uid35_bh7_uid36_In0: (c0, 1.100000ns)
signal Compressor_14_3_Freq200_uid35_bh7_uid36_In1 :  std_logic_vector(0 downto 0);
   -- timing of Compressor_14_3_Freq200_uid35_bh7_uid36_In1: (c0, 1.100000ns)
signal Compressor_14_3_Freq200_uid35_bh7_uid36_Out0 :  std_logic_vector(2 downto 0);
   -- timing of Compressor_14_3_Freq200_uid35_bh7_uid36_Out0: (c0, 1.650000ns)
signal bh7_w14_3 :  std_logic;
   -- timing of bh7_w14_3: (c0, 1.650000ns)
signal bh7_w15_1 :  std_logic;
   -- timing of bh7_w15_1: (c0, 1.650000ns)
signal bh7_w16_1 :  std_logic;
   -- timing of bh7_w16_1: (c0, 1.650000ns)
signal Compressor_14_3_Freq200_uid35_bh7_uid36_Out0_copy37 :  std_logic_vector(2 downto 0);
   -- timing of Compressor_14_3_Freq200_uid35_bh7_uid36_Out0_copy37: (c0, 1.100000ns)
signal tmp_bitheapResult_bh7_0 :  std_logic_vector(0 downto 0);
   -- timing of tmp_bitheapResult_bh7_0: (c0, 1.700000ns)
signal bitheapFinalAdd_bh7_In0 :  std_logic_vector(18 downto 0);
   -- timing of bitheapFinalAdd_bh7_In0: (c0, 1.700000ns)
signal bitheapFinalAdd_bh7_In1 :  std_logic_vector(18 downto 0);
   -- timing of bitheapFinalAdd_bh7_In1: (c0, 1.700000ns)
signal bitheapFinalAdd_bh7_Cin :  std_logic;
   -- timing of bitheapFinalAdd_bh7_Cin: (c0, 0.000000ns)
signal bitheapFinalAdd_bh7_Out :  std_logic_vector(18 downto 0);
   -- timing of bitheapFinalAdd_bh7_Out: (c0, 2.880000ns)
signal bitheapResult_bh7 :  std_logic_vector(19 downto 0);
   -- timing of bitheapResult_bh7: (c0, 2.880000ns)
signal OutRes :  std_logic_vector(19 downto 0);
   -- timing of OutRes: (c0, 2.880000ns)
begin
-- This operator multiplies by pi
   FixRealKCM_Freq200_uid6_A0 <= X(15 downto 11);-- input address  m=-13  l=-17
   FixRealKCM_Freq200_uid6_Table0: FixRealKCM_Freq200_uid6_T0_Freq200_uid9
      port map ( X => FixRealKCM_Freq200_uid6_A0,
                 Y => FixRealKCM_Freq200_uid6_T0_copy10);
   FixRealKCM_Freq200_uid6_T0 <= FixRealKCM_Freq200_uid6_T0_copy10; -- output copy to hold a pipeline register if needed
   bh7_w0_0 <= FixRealKCM_Freq200_uid6_T0(0);
   bh7_w1_0 <= FixRealKCM_Freq200_uid6_T0(1);
   bh7_w2_0 <= FixRealKCM_Freq200_uid6_T0(2);
   bh7_w3_0 <= FixRealKCM_Freq200_uid6_T0(3);
   bh7_w4_0 <= FixRealKCM_Freq200_uid6_T0(4);
   bh7_w5_0 <= FixRealKCM_Freq200_uid6_T0(5);
   bh7_w6_0 <= FixRealKCM_Freq200_uid6_T0(6);
   bh7_w7_0 <= FixRealKCM_Freq200_uid6_T0(7);
   bh7_w8_0 <= FixRealKCM_Freq200_uid6_T0(8);
   bh7_w9_0 <= FixRealKCM_Freq200_uid6_T0(9);
   bh7_w10_0 <= FixRealKCM_Freq200_uid6_T0(10);
   bh7_w11_0 <= FixRealKCM_Freq200_uid6_T0(11);
   bh7_w12_0 <= FixRealKCM_Freq200_uid6_T0(12);
   bh7_w13_0 <= FixRealKCM_Freq200_uid6_T0(13);
   bh7_w14_0 <= FixRealKCM_Freq200_uid6_T0(14);
   bh7_w15_0 <= FixRealKCM_Freq200_uid6_T0(15);
   bh7_w16_0 <= FixRealKCM_Freq200_uid6_T0(16);
   bh7_w17_0 <= FixRealKCM_Freq200_uid6_T0(17);
   bh7_w18_0 <= FixRealKCM_Freq200_uid6_T0(18);
   bh7_w19_0 <= FixRealKCM_Freq200_uid6_T0(19);
   FixRealKCM_Freq200_uid6_A1 <= X(10 downto 6);-- input address  m=-18  l=-22
   FixRealKCM_Freq200_uid6_Table1: FixRealKCM_Freq200_uid6_T1_Freq200_uid12
      port map ( X => FixRealKCM_Freq200_uid6_A1,
                 Y => FixRealKCM_Freq200_uid6_T1_copy13);
   FixRealKCM_Freq200_uid6_T1 <= FixRealKCM_Freq200_uid6_T1_copy13; -- output copy to hold a pipeline register if needed
   bh7_w0_1 <= FixRealKCM_Freq200_uid6_T1(0);
   bh7_w1_1 <= FixRealKCM_Freq200_uid6_T1(1);
   bh7_w2_1 <= FixRealKCM_Freq200_uid6_T1(2);
   bh7_w3_1 <= FixRealKCM_Freq200_uid6_T1(3);
   bh7_w4_1 <= FixRealKCM_Freq200_uid6_T1(4);
   bh7_w5_1 <= FixRealKCM_Freq200_uid6_T1(5);
   bh7_w6_1 <= FixRealKCM_Freq200_uid6_T1(6);
   bh7_w7_1 <= FixRealKCM_Freq200_uid6_T1(7);
   bh7_w8_1 <= FixRealKCM_Freq200_uid6_T1(8);
   bh7_w9_1 <= FixRealKCM_Freq200_uid6_T1(9);
   bh7_w10_1 <= FixRealKCM_Freq200_uid6_T1(10);
   bh7_w11_1 <= FixRealKCM_Freq200_uid6_T1(11);
   bh7_w12_1 <= FixRealKCM_Freq200_uid6_T1(12);
   bh7_w13_1 <= FixRealKCM_Freq200_uid6_T1(13);
   bh7_w14_1 <= FixRealKCM_Freq200_uid6_T1(14);
   FixRealKCM_Freq200_uid6_A2 <= X(5 downto 0);-- input address  m=-23  l=-28
   FixRealKCM_Freq200_uid6_Table2: FixRealKCM_Freq200_uid6_T2_Freq200_uid15
      port map ( X => FixRealKCM_Freq200_uid6_A2,
                 Y => FixRealKCM_Freq200_uid6_T2_copy16);
   FixRealKCM_Freq200_uid6_T2 <= FixRealKCM_Freq200_uid6_T2_copy16; -- output copy to hold a pipeline register if needed
   bh7_w0_2 <= FixRealKCM_Freq200_uid6_T2(0);
   bh7_w1_2 <= FixRealKCM_Freq200_uid6_T2(1);
   bh7_w2_2 <= FixRealKCM_Freq200_uid6_T2(2);
   bh7_w3_2 <= FixRealKCM_Freq200_uid6_T2(3);
   bh7_w4_2 <= FixRealKCM_Freq200_uid6_T2(4);
   bh7_w5_2 <= FixRealKCM_Freq200_uid6_T2(5);
   bh7_w6_2 <= FixRealKCM_Freq200_uid6_T2(6);
   bh7_w7_2 <= FixRealKCM_Freq200_uid6_T2(7);
   bh7_w8_2 <= FixRealKCM_Freq200_uid6_T2(8);
   bh7_w9_2 <= FixRealKCM_Freq200_uid6_T2(9);

   -- Adding the constant bits 
      -- All the constant bits are zero, nothing to add


   Compressor_23_3_Freq200_uid19_bh7_uid20_In0 <= "" & bh7_w0_1 & bh7_w0_0 & bh7_w0_2;
   Compressor_23_3_Freq200_uid19_bh7_uid20_In1 <= "" & bh7_w1_1 & bh7_w1_0;
   bh7_w0_3 <= Compressor_23_3_Freq200_uid19_bh7_uid20_Out0(0);
   bh7_w1_3 <= Compressor_23_3_Freq200_uid19_bh7_uid20_Out0(1);
   bh7_w2_3 <= Compressor_23_3_Freq200_uid19_bh7_uid20_Out0(2);
   Compressor_23_3_Freq200_uid19_uid20: Compressor_23_3_Freq200_uid19
      port map ( X0 => Compressor_23_3_Freq200_uid19_bh7_uid20_In0,
                 X1 => Compressor_23_3_Freq200_uid19_bh7_uid20_In1,
                 R => Compressor_23_3_Freq200_uid19_bh7_uid20_Out0_copy21);
   Compressor_23_3_Freq200_uid19_bh7_uid20_Out0 <= Compressor_23_3_Freq200_uid19_bh7_uid20_Out0_copy21; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq200_uid19_bh7_uid22_In0 <= "" & bh7_w2_1 & bh7_w2_0 & bh7_w2_2;
   Compressor_23_3_Freq200_uid19_bh7_uid22_In1 <= "" & bh7_w3_1 & bh7_w3_0;
   bh7_w2_4 <= Compressor_23_3_Freq200_uid19_bh7_uid22_Out0(0);
   bh7_w3_3 <= Compressor_23_3_Freq200_uid19_bh7_uid22_Out0(1);
   bh7_w4_3 <= Compressor_23_3_Freq200_uid19_bh7_uid22_Out0(2);
   Compressor_23_3_Freq200_uid19_uid22: Compressor_23_3_Freq200_uid19
      port map ( X0 => Compressor_23_3_Freq200_uid19_bh7_uid22_In0,
                 X1 => Compressor_23_3_Freq200_uid19_bh7_uid22_In1,
                 R => Compressor_23_3_Freq200_uid19_bh7_uid22_Out0_copy23);
   Compressor_23_3_Freq200_uid19_bh7_uid22_Out0 <= Compressor_23_3_Freq200_uid19_bh7_uid22_Out0_copy23; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq200_uid19_bh7_uid24_In0 <= "" & bh7_w4_1 & bh7_w4_0 & bh7_w4_2;
   Compressor_23_3_Freq200_uid19_bh7_uid24_In1 <= "" & bh7_w5_1 & bh7_w5_0;
   bh7_w4_4 <= Compressor_23_3_Freq200_uid19_bh7_uid24_Out0(0);
   bh7_w5_3 <= Compressor_23_3_Freq200_uid19_bh7_uid24_Out0(1);
   bh7_w6_3 <= Compressor_23_3_Freq200_uid19_bh7_uid24_Out0(2);
   Compressor_23_3_Freq200_uid19_uid24: Compressor_23_3_Freq200_uid19
      port map ( X0 => Compressor_23_3_Freq200_uid19_bh7_uid24_In0,
                 X1 => Compressor_23_3_Freq200_uid19_bh7_uid24_In1,
                 R => Compressor_23_3_Freq200_uid19_bh7_uid24_Out0_copy25);
   Compressor_23_3_Freq200_uid19_bh7_uid24_Out0 <= Compressor_23_3_Freq200_uid19_bh7_uid24_Out0_copy25; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq200_uid19_bh7_uid26_In0 <= "" & bh7_w6_1 & bh7_w6_0 & bh7_w6_2;
   Compressor_23_3_Freq200_uid19_bh7_uid26_In1 <= "" & bh7_w7_1 & bh7_w7_0;
   bh7_w6_4 <= Compressor_23_3_Freq200_uid19_bh7_uid26_Out0(0);
   bh7_w7_3 <= Compressor_23_3_Freq200_uid19_bh7_uid26_Out0(1);
   bh7_w8_3 <= Compressor_23_3_Freq200_uid19_bh7_uid26_Out0(2);
   Compressor_23_3_Freq200_uid19_uid26: Compressor_23_3_Freq200_uid19
      port map ( X0 => Compressor_23_3_Freq200_uid19_bh7_uid26_In0,
                 X1 => Compressor_23_3_Freq200_uid19_bh7_uid26_In1,
                 R => Compressor_23_3_Freq200_uid19_bh7_uid26_Out0_copy27);
   Compressor_23_3_Freq200_uid19_bh7_uid26_Out0 <= Compressor_23_3_Freq200_uid19_bh7_uid26_Out0_copy27; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq200_uid19_bh7_uid28_In0 <= "" & bh7_w8_1 & bh7_w8_0 & bh7_w8_2;
   Compressor_23_3_Freq200_uid19_bh7_uid28_In1 <= "" & bh7_w9_1 & bh7_w9_0;
   bh7_w8_4 <= Compressor_23_3_Freq200_uid19_bh7_uid28_Out0(0);
   bh7_w9_3 <= Compressor_23_3_Freq200_uid19_bh7_uid28_Out0(1);
   bh7_w10_2 <= Compressor_23_3_Freq200_uid19_bh7_uid28_Out0(2);
   Compressor_23_3_Freq200_uid19_uid28: Compressor_23_3_Freq200_uid19
      port map ( X0 => Compressor_23_3_Freq200_uid19_bh7_uid28_In0,
                 X1 => Compressor_23_3_Freq200_uid19_bh7_uid28_In1,
                 R => Compressor_23_3_Freq200_uid19_bh7_uid28_Out0_copy29);
   Compressor_23_3_Freq200_uid19_bh7_uid28_Out0 <= Compressor_23_3_Freq200_uid19_bh7_uid28_Out0_copy29; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq200_uid19_bh7_uid30_In0 <= "" & bh7_w10_1 & bh7_w10_0 & "0";
   Compressor_23_3_Freq200_uid19_bh7_uid30_In1 <= "" & bh7_w11_1 & bh7_w11_0;
   bh7_w10_3 <= Compressor_23_3_Freq200_uid19_bh7_uid30_Out0(0);
   bh7_w11_2 <= Compressor_23_3_Freq200_uid19_bh7_uid30_Out0(1);
   bh7_w12_2 <= Compressor_23_3_Freq200_uid19_bh7_uid30_Out0(2);
   Compressor_23_3_Freq200_uid19_uid30: Compressor_23_3_Freq200_uid19
      port map ( X0 => Compressor_23_3_Freq200_uid19_bh7_uid30_In0,
                 X1 => Compressor_23_3_Freq200_uid19_bh7_uid30_In1,
                 R => Compressor_23_3_Freq200_uid19_bh7_uid30_Out0_copy31);
   Compressor_23_3_Freq200_uid19_bh7_uid30_Out0 <= Compressor_23_3_Freq200_uid19_bh7_uid30_Out0_copy31; -- output copy to hold a pipeline register if needed


   Compressor_23_3_Freq200_uid19_bh7_uid32_In0 <= "" & bh7_w12_1 & bh7_w12_0 & "0";
   Compressor_23_3_Freq200_uid19_bh7_uid32_In1 <= "" & bh7_w13_1 & bh7_w13_0;
   bh7_w12_3 <= Compressor_23_3_Freq200_uid19_bh7_uid32_Out0(0);
   bh7_w13_2 <= Compressor_23_3_Freq200_uid19_bh7_uid32_Out0(1);
   bh7_w14_2 <= Compressor_23_3_Freq200_uid19_bh7_uid32_Out0(2);
   Compressor_23_3_Freq200_uid19_uid32: Compressor_23_3_Freq200_uid19
      port map ( X0 => Compressor_23_3_Freq200_uid19_bh7_uid32_In0,
                 X1 => Compressor_23_3_Freq200_uid19_bh7_uid32_In1,
                 R => Compressor_23_3_Freq200_uid19_bh7_uid32_Out0_copy33);
   Compressor_23_3_Freq200_uid19_bh7_uid32_Out0 <= Compressor_23_3_Freq200_uid19_bh7_uid32_Out0_copy33; -- output copy to hold a pipeline register if needed


   Compressor_14_3_Freq200_uid35_bh7_uid36_In0 <= "" & bh7_w14_1 & bh7_w14_0 & "0" & "0";
   Compressor_14_3_Freq200_uid35_bh7_uid36_In1 <= "" & bh7_w15_0;
   bh7_w14_3 <= Compressor_14_3_Freq200_uid35_bh7_uid36_Out0(0);
   bh7_w15_1 <= Compressor_14_3_Freq200_uid35_bh7_uid36_Out0(1);
   bh7_w16_1 <= Compressor_14_3_Freq200_uid35_bh7_uid36_Out0(2);
   Compressor_14_3_Freq200_uid35_uid36: Compressor_14_3_Freq200_uid35
      port map ( X0 => Compressor_14_3_Freq200_uid35_bh7_uid36_In0,
                 X1 => Compressor_14_3_Freq200_uid35_bh7_uid36_In1,
                 R => Compressor_14_3_Freq200_uid35_bh7_uid36_Out0_copy37);
   Compressor_14_3_Freq200_uid35_bh7_uid36_Out0 <= Compressor_14_3_Freq200_uid35_bh7_uid36_Out0_copy37; -- output copy to hold a pipeline register if needed

   tmp_bitheapResult_bh7_0(0) <= bh7_w0_3;

   bitheapFinalAdd_bh7_In0 <= "" & bh7_w19_0 & bh7_w18_0 & bh7_w17_0 & bh7_w16_0 & bh7_w15_1 & bh7_w14_3 & bh7_w13_2 & bh7_w12_3 & bh7_w11_2 & bh7_w10_3 & bh7_w9_2 & bh7_w8_4 & bh7_w7_2 & bh7_w6_4 & bh7_w5_2 & bh7_w4_4 & bh7_w3_2 & bh7_w2_4 & bh7_w1_2;
   bitheapFinalAdd_bh7_In1 <= "0" & "0" & "0" & bh7_w16_1 & "0" & bh7_w14_2 & "0" & bh7_w12_2 & "0" & bh7_w10_2 & bh7_w9_3 & bh7_w8_3 & bh7_w7_3 & bh7_w6_3 & bh7_w5_3 & bh7_w4_3 & bh7_w3_3 & bh7_w2_3 & bh7_w1_3;
   bitheapFinalAdd_bh7_Cin <= '0';

   bitheapFinalAdd_bh7: IntAdder_19_Freq200_uid39
      port map ( clk  => clk,
                 rst  => rst,
                 Cin => bitheapFinalAdd_bh7_Cin,
                 X => bitheapFinalAdd_bh7_In0,
                 Y => bitheapFinalAdd_bh7_In1,
                 R => bitheapFinalAdd_bh7_Out);
   bitheapResult_bh7 <= bitheapFinalAdd_bh7_Out(18 downto 0) & tmp_bitheapResult_bh7_0;
   OutRes <= bitheapResult_bh7(19 downto 0);
   R <= OutRes(19 downto 2);
end architecture;

--------------------------------------------------------------------------------
--                                FixSinCos_24
--                    (FixSinCosPoly_LSBm24_Freq200_uid2)
-- VHDL generated for DummyFPGA @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Antoine Martinet, Guillaume Sergent, (2013-2019)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: S C
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: S: (c2, 3.029062ns)C: (c2, 3.029062ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixSinCos_24 is
    port (clk, rst : in std_logic;
          X : in  std_logic_vector(24 downto 0);
          S : out  std_logic_vector(24 downto 0);
          C : out  std_logic_vector(24 downto 0)   );
end entity;

architecture arch of FixSinCos_24 is
   component SinCosTable_Freq200_uid4 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(9 downto 0);
             Y : out  std_logic_vector(55 downto 0)   );
   end component;

   component FixRealKCM_Freq200_uid6 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(15 downto 0);
             R : out  std_logic_vector(17 downto 0)   );
   end component;

   component FixFunctionByTable_Freq200_uid41 is
      port ( X : in  std_logic_vector(6 downto 0);
             Y : out  std_logic_vector(6 downto 0)   );
   end component;

signal X_sgn, X_sgn_d1, X_sgn_d2 :  std_logic;
   -- timing of X_sgn: (c0, 0.000000ns)
signal Q :  std_logic;
   -- timing of Q: (c0, 0.000000ns)
signal O :  std_logic;
   -- timing of O: (c0, 0.000000ns)
signal Y :  std_logic_vector(21 downto 0);
   -- timing of Y: (c0, 0.000000ns)
signal Yneg :  std_logic_vector(25 downto 0);
   -- timing of Yneg: (c0, 0.550000ns)
signal A :  std_logic_vector(9 downto 0);
   -- timing of A: (c0, 0.550000ns)
signal Y_red :  std_logic_vector(15 downto 0);
   -- timing of Y_red: (c0, 0.550000ns)
signal SinCosA :  std_logic_vector(55 downto 0);
   -- timing of SinCosA: (c1, 2.789062ns)
signal SinPiA, SinPiA_d1 :  std_logic_vector(27 downto 0);
   -- timing of SinPiA: (c1, 2.789062ns)
signal CosPiA, CosPiA_d1 :  std_logic_vector(27 downto 0);
   -- timing of CosPiA: (c1, 2.789062ns)
signal Z, Z_d1, Z_d2 :  std_logic_vector(17 downto 0);
   -- timing of Z: (c0, 2.880000ns)
signal Z_trunc_for_square :  std_logic_vector(6 downto 0);
   -- timing of Z_trunc_for_square: (c0, 2.880000ns)
signal Z2o2_w :  std_logic_vector(6 downto 0);
   -- timing of Z2o2_w: (c0, 3.430000ns)
signal Z2o2_w_copy42 :  std_logic_vector(6 downto 0);
   -- timing of Z2o2_w_copy42: (c0, 2.880000ns)
signal Z2o2, Z2o2_d1, Z2o2_d2 :  std_logic_vector(6 downto 0);
   -- timing of Z2o2: (c0, 3.430000ns)
signal CosPiA_trunc_to_z2o2, CosPiA_trunc_to_z2o2_d1 :  std_logic_vector(6 downto 0);
   -- timing of CosPiA_trunc_to_z2o2: (c1, 2.789062ns)
signal Z2o2CosPiA :  std_logic_vector(13 downto 0);
   -- timing of Z2o2CosPiA: (c2, 0.489062ns)
signal Z2o2CosPiA_aligned :  std_logic_vector(27 downto 0);
   -- timing of Z2o2CosPiA_aligned: (c2, 0.489062ns)
signal CosPiACosZ :  std_logic_vector(27 downto 0);
   -- timing of CosPiACosZ: (c2, 1.759062ns)
signal SinPiA_trunc_to_z2o2, SinPiA_trunc_to_z2o2_d1 :  std_logic_vector(6 downto 0);
   -- timing of SinPiA_trunc_to_z2o2: (c1, 2.789062ns)
signal Z2o2SinPiA :  std_logic_vector(13 downto 0);
   -- timing of Z2o2SinPiA: (c2, 0.489062ns)
signal Z2o2SinPiA_aligned :  std_logic_vector(27 downto 0);
   -- timing of Z2o2SinPiA_aligned: (c2, 0.489062ns)
signal SinPiACosZ :  std_logic_vector(27 downto 0);
   -- timing of SinPiACosZ: (c2, 1.759062ns)
signal CosPiAZ :  std_logic_vector(45 downto 0);
   -- timing of CosPiAZ: (c2, 0.489062ns)
signal CosPiASinZ :  std_logic_vector(27 downto 0);
   -- timing of CosPiASinZ: (c2, 0.489062ns)
signal SinPiAZ :  std_logic_vector(45 downto 0);
   -- timing of SinPiAZ: (c2, 0.489062ns)
signal SinPiASinZ :  std_logic_vector(27 downto 0);
   -- timing of SinPiASinZ: (c2, 0.489062ns)
signal PreSinX :  std_logic_vector(27 downto 0);
   -- timing of PreSinX: (c2, 3.029062ns)
signal PreCosX :  std_logic_vector(27 downto 0);
   -- timing of PreCosX: (c2, 3.029062ns)
signal C_out :  std_logic_vector(23 downto 0);
   -- timing of C_out: (c2, 3.029062ns)
signal S_out :  std_logic_vector(23 downto 0);
   -- timing of S_out: (c2, 3.029062ns)
signal C_sgn, C_sgn_d1, C_sgn_d2 :  std_logic;
   -- timing of C_sgn: (c0, 0.000000ns)
signal Exch, Exch_d1, Exch_d2 :  std_logic;
   -- timing of Exch: (c0, 0.000000ns)
signal S_wo_sgn :  std_logic_vector(23 downto 0);
   -- timing of S_wo_sgn: (c2, 3.029062ns)
signal C_wo_sgn :  std_logic_vector(23 downto 0);
   -- timing of C_wo_sgn: (c2, 3.029062ns)
signal S_wo_sgn_ext :  std_logic_vector(24 downto 0);
   -- timing of S_wo_sgn_ext: (c2, 3.029062ns)
signal C_wo_sgn_ext :  std_logic_vector(24 downto 0);
   -- timing of C_wo_sgn_ext: (c2, 3.029062ns)
signal S_wo_sgn_neg :  std_logic_vector(24 downto 0);
   -- timing of S_wo_sgn_neg: (c2, 3.029062ns)
signal C_wo_sgn_neg :  std_logic_vector(24 downto 0);
   -- timing of C_wo_sgn_neg: (c2, 3.029062ns)
begin
   process(clk, rst)
      begin
         if rst = '1' then
            X_sgn_d1 <=  '0';
            X_sgn_d2 <=  '0';
            SinPiA_d1 <=  (others => '0');
            CosPiA_d1 <=  (others => '0');
            Z_d1 <=  (others => '0');
            Z_d2 <=  (others => '0');
            Z2o2_d1 <=  (others => '0');
            Z2o2_d2 <=  (others => '0');
            CosPiA_trunc_to_z2o2_d1 <=  (others => '0');
            SinPiA_trunc_to_z2o2_d1 <=  (others => '0');
            C_sgn_d1 <=  '0';
            C_sgn_d2 <=  '0';
            Exch_d1 <=  '0';
            Exch_d2 <=  '0';
         elsif clk'event and clk = '1' then
            X_sgn_d1 <=  X_sgn;
            X_sgn_d2 <=  X_sgn_d1;
            SinPiA_d1 <=  SinPiA;
            CosPiA_d1 <=  CosPiA;
            Z_d1 <=  Z;
            Z_d2 <=  Z_d1;
            Z2o2_d1 <=  Z2o2;
            Z2o2_d2 <=  Z2o2_d1;
            CosPiA_trunc_to_z2o2_d1 <=  CosPiA_trunc_to_z2o2;
            SinPiA_trunc_to_z2o2_d1 <=  SinPiA_trunc_to_z2o2;
            C_sgn_d1 <=  C_sgn;
            C_sgn_d2 <=  C_sgn_d1;
            Exch_d1 <=  Exch;
            Exch_d2 <=  Exch_d1;
         end if;
      end process;
   -- The argument is reduced into (0,1/4)
   X_sgn <= X(24);  -- sign
   Q <= X(23);  -- quadrant
   O <= X(22);  -- octant
   Y <= X (21 downto 0);
   -- Computing .25-Y :  we do a logic NOT, at a cost of 1 ulp
   Yneg <= ((not Y) & "1111") when O='1' else (Y & "0000");
   A <= Yneg (25 downto 16);
   Y_red <= Yneg(15 downto 0);
   SinCosTable: SinCosTable_Freq200_uid4
      port map ( clk  => clk,
                 rst  => rst,
                 X => A,
                 Y => SinCosA);
   SinPiA <= SinCosA(55 downto 28);
   CosPiA <= SinCosA(27 downto 0);
   MultByPi: FixRealKCM_Freq200_uid6
      port map ( clk  => clk,
                 rst  => rst,
                 X => Y_red,
                 R => Z);
   Z_trunc_for_square<= Z (17 downto 11);
   ZSquarer: FixFunctionByTable_Freq200_uid41
      port map ( X => Z_trunc_for_square,
                 Y => Z2o2_w_copy42);
   Z2o2_w <= Z2o2_w_copy42; -- output copy to hold a pipeline register if needed
   Z2o2 <= Z2o2_w(6 downto 0); -- get rid of the possible constant 0
   CosPiA_trunc_to_z2o2 <= CosPiA(27 downto 21);
   Z2o2CosPiA <=  CosPiA_trunc_to_z2o2_d1 * Z2o2_d2;
   Z2o2CosPiA_aligned <= "000000000000000000000" & Z2o2CosPiA(13 downto 7);
   CosPiACosZ<= CosPiA_d1 - Z2o2CosPiA_aligned;
   SinPiA_trunc_to_z2o2 <= SinPiA(27 downto 21);
   Z2o2SinPiA <=  SinPiA_trunc_to_z2o2_d1 * Z2o2_d2;
   Z2o2SinPiA_aligned <= "000000000000000000000" & Z2o2SinPiA(13 downto 7);
   SinPiACosZ<= SinPiA_d1 - Z2o2SinPiA_aligned;
   CosPiAZ <= CosPiA_d1*Z_d2;  -- TODO check it fits DSP
   CosPiASinZ <= "0000000000" & CosPiAZ(45 downto 28);
   SinPiAZ <= SinPiA_d1*Z_d2;  -- TODO check it fits DSP
   SinPiASinZ <= "0000000000" & SinPiAZ(45 downto 28);
   PreSinX <= SinPiACosZ + CosPiASinZ;
   PreCosX <= CosPiACosZ - SinPiASinZ;
   C_out <= PreCosX(27 downto 4);
   S_out <= PreSinX(27 downto 4);
   -- --- Final reconstruction of both sine and cosine ---
   C_sgn <= X_sgn xor Q;
   Exch <= Q xor O;
   S_wo_sgn <= C_out when Exch_d2 = '1' else S_out;
   C_wo_sgn <= S_out when Exch_d2 = '1' else C_out;
   S_wo_sgn_ext <= '0' & S_wo_sgn;
   C_wo_sgn_ext <= '0' & C_wo_sgn;
   S_wo_sgn_neg <= (not S_wo_sgn_ext) + 1;
   C_wo_sgn_neg <= (not C_wo_sgn_ext) + 1;
   S <= S_wo_sgn_ext when X_sgn_d2 = '0' else S_wo_sgn_neg;
   C <= C_wo_sgn_ext when C_sgn_d2 = '0' else C_wo_sgn_neg;
end architecture;

