--------------------------------------------------------------------------------
--                          SinCosTable_Freq200_uid4
-- VHDL generated for DummyFPGA @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007-2022)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: Y
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: Y: (c1, 2.239062ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity SinCosTable_Freq200_uid4 is
    port (clk, rst : in std_logic;
          X : in  std_logic_vector(9 downto 0);
          Y : out  std_logic_vector(21 downto 0)   );
end entity;

architecture arch of SinCosTable_Freq200_uid4 is
signal Y0, Y0_d1 :  std_logic_vector(21 downto 0);
   -- timing of Y0: (c0, 2.000000ns)
signal Y1 :  std_logic_vector(21 downto 0);
   -- timing of Y1: (c1, 2.239062ns)
begin
   process(clk, rst)
      begin
         if rst = '1' then
            Y0_d1 <=  (others => '0');
         elsif clk'event and clk = '1' then
            Y0_d1 <=  Y0;
         end if;
      end process;
   with X  select  Y0 <= 
      "0000000000011111111111" when "0000000000",
      "0000000001111111111111" when "0000000001",
      "0000000011011111111111" when "0000000010",
      "0000000100111111111111" when "0000000011",
      "0000000110111111111111" when "0000000100",
      "0000001000011111111111" when "0000000101",
      "0000001001111111111111" when "0000000110",
      "0000001011011111111111" when "0000000111",
      "0000001100111111111111" when "0000001000",
      "0000001110011111111111" when "0000001001",
      "0000001111111111111111" when "0000001010",
      "0000010001111111111111" when "0000001011",
      "0000010011011111111111" when "0000001100",
      "0000010100111111111111" when "0000001101",
      "0000010110011111111111" when "0000001110",
      "0000010111111111111110" when "0000001111",
      "0000011001011111111110" when "0000010000",
      "0000011010111111111110" when "0000010001",
      "0000011100111111111110" when "0000010010",
      "0000011110011111111110" when "0000010011",
      "0000011111111111111110" when "0000010100",
      "0000100001011111111110" when "0000010101",
      "0000100010111111111110" when "0000010110",
      "0000100100011111111110" when "0000010111",
      "0000100101111111111110" when "0000011000",
      "0000100111011111111101" when "0000011001",
      "0000101001011111111101" when "0000011010",
      "0000101010111111111101" when "0000011011",
      "0000101100011111111101" when "0000011100",
      "0000101101111111111101" when "0000011101",
      "0000101111011111111101" when "0000011110",
      "0000110000111111111101" when "0000011111",
      "0000110010011111111101" when "0000100000",
      "0000110100011111111100" when "0000100001",
      "0000110101111111111100" when "0000100010",
      "0000110111011111111100" when "0000100011",
      "0000111000111111111100" when "0000100100",
      "0000111010011111111100" when "0000100101",
      "0000111011111111111100" when "0000100110",
      "0000111101011111111011" when "0000100111",
      "0000111111011111111011" when "0000101000",
      "0001000000111111111011" when "0000101001",
      "0001000010011111111011" when "0000101010",
      "0001000011111111111011" when "0000101011",
      "0001000101011111111010" when "0000101100",
      "0001000110111111111010" when "0000101101",
      "0001001000011111111010" when "0000101110",
      "0001001001111111111010" when "0000101111",
      "0001001011111111111001" when "0000110000",
      "0001001101011111111001" when "0000110001",
      "0001001110111111111001" when "0000110010",
      "0001010000011111111001" when "0000110011",
      "0001010001111111111000" when "0000110100",
      "0001010011011111111000" when "0000110101",
      "0001010100111111111000" when "0000110110",
      "0001010110011111111000" when "0000110111",
      "0001011000011111110111" when "0000111000",
      "0001011001111111110111" when "0000111001",
      "0001011011011111110111" when "0000111010",
      "0001011100111111110111" when "0000111011",
      "0001011110011111110110" when "0000111100",
      "0001011111111111110110" when "0000111101",
      "0001100001011111110110" when "0000111110",
      "0001100011011111110101" when "0000111111",
      "0001100100111111110101" when "0001000000",
      "0001100110011111110101" when "0001000001",
      "0001100111111111110101" when "0001000010",
      "0001101001011111110100" when "0001000011",
      "0001101010111111110100" when "0001000100",
      "0001101100011111110100" when "0001000101",
      "0001101101111111110011" when "0001000110",
      "0001101111111111110011" when "0001000111",
      "0001110001011111110011" when "0001001000",
      "0001110010111111110010" when "0001001001",
      "0001110100011111110010" when "0001001010",
      "0001110101111111110001" when "0001001011",
      "0001110111011111110001" when "0001001100",
      "0001111000111111110001" when "0001001101",
      "0001111010011111110000" when "0001001110",
      "0001111011111111110000" when "0001001111",
      "0001111101111111110000" when "0001010000",
      "0001111111011111101111" when "0001010001",
      "0010000000111111101111" when "0001010010",
      "0010000010011111101110" when "0001010011",
      "0010000011111111101110" when "0001010100",
      "0010000101011111101110" when "0001010101",
      "0010000110111111101101" when "0001010110",
      "0010001000011111101101" when "0001010111",
      "0010001001111111101100" when "0001011000",
      "0010001011111111101100" when "0001011001",
      "0010001101011111101100" when "0001011010",
      "0010001110111111101011" when "0001011011",
      "0010010000011111101011" when "0001011100",
      "0010010001111111101010" when "0001011101",
      "0010010011011111101010" when "0001011110",
      "0010010100111111101001" when "0001011111",
      "0010010110011111101001" when "0001100000",
      "0010010111111111101000" when "0001100001",
      "0010011001111111101000" when "0001100010",
      "0010011011011111100111" when "0001100011",
      "0010011100111111100111" when "0001100100",
      "0010011110011111100110" when "0001100101",
      "0010011111111111100110" when "0001100110",
      "0010100001011111100110" when "0001100111",
      "0010100010111111100101" when "0001101000",
      "0010100100011111100101" when "0001101001",
      "0010100101111111100100" when "0001101010",
      "0010100111011111100011" when "0001101011",
      "0010101001011111100011" when "0001101100",
      "0010101010111111100010" when "0001101101",
      "0010101100011111100010" when "0001101110",
      "0010101101111111100001" when "0001101111",
      "0010101111011111100001" when "0001110000",
      "0010110000111111100000" when "0001110001",
      "0010110010011111100000" when "0001110010",
      "0010110011111111011111" when "0001110011",
      "0010110101011111011111" when "0001110100",
      "0010110110111111011110" when "0001110101",
      "0010111000111111011110" when "0001110110",
      "0010111010011111011101" when "0001110111",
      "0010111011111111011100" when "0001111000",
      "0010111101011111011100" when "0001111001",
      "0010111110111111011011" when "0001111010",
      "0011000000011111011011" when "0001111011",
      "0011000001111111011010" when "0001111100",
      "0011000011011111011001" when "0001111101",
      "0011000100111111011001" when "0001111110",
      "0011000110011111011000" when "0001111111",
      "0011000111111111011000" when "0010000000",
      "0011001001011111010111" when "0010000001",
      "0011001011011111010110" when "0010000010",
      "0011001100111111010110" when "0010000011",
      "0011001110011111010101" when "0010000100",
      "0011001111111111010101" when "0010000101",
      "0011010001011111010100" when "0010000110",
      "0011010010111111010011" when "0010000111",
      "0011010100011111010011" when "0010001000",
      "0011010101111111010010" when "0010001001",
      "0011010111011111010001" when "0010001010",
      "0011011000111111010001" when "0010001011",
      "0011011010011111010000" when "0010001100",
      "0011011011111111001111" when "0010001101",
      "0011011101011111001111" when "0010001110",
      "0011011110111111001110" when "0010001111",
      "0011100000111111001101" when "0010010000",
      "0011100010011111001101" when "0010010001",
      "0011100011111111001100" when "0010010010",
      "0011100101011111001011" when "0010010011",
      "0011100110111111001010" when "0010010100",
      "0011101000011111001010" when "0010010101",
      "0011101001111111001001" when "0010010110",
      "0011101011011111001000" when "0010010111",
      "0011101100111111001000" when "0010011000",
      "0011101110011111000111" when "0010011001",
      "0011101111111111000110" when "0010011010",
      "0011110001011111000101" when "0010011011",
      "0011110010111111000101" when "0010011100",
      "0011110100011111000100" when "0010011101",
      "0011110101111111000011" when "0010011110",
      "0011110111011111000010" when "0010011111",
      "0011111000111111000010" when "0010100000",
      "0011111010011111000001" when "0010100001",
      "0011111011111111000000" when "0010100010",
      "0011111101111110111111" when "0010100011",
      "0011111111011110111111" when "0010100100",
      "0100000000111110111110" when "0010100101",
      "0100000010011110111101" when "0010100110",
      "0100000011111110111100" when "0010100111",
      "0100000101011110111011" when "0010101000",
      "0100000110111110111011" when "0010101001",
      "0100001000011110111010" when "0010101010",
      "0100001001111110111001" when "0010101011",
      "0100001011011110111000" when "0010101100",
      "0100001100111110110111" when "0010101101",
      "0100001110011110110111" when "0010101110",
      "0100001111111110110110" when "0010101111",
      "0100010001011110110101" when "0010110000",
      "0100010010111110110100" when "0010110001",
      "0100010100011110110011" when "0010110010",
      "0100010101111110110010" when "0010110011",
      "0100010111011110110001" when "0010110100",
      "0100011000111110110001" when "0010110101",
      "0100011010011110110000" when "0010110110",
      "0100011011111110101111" when "0010110111",
      "0100011101011110101110" when "0010111000",
      "0100011110111110101101" when "0010111001",
      "0100100000011110101100" when "0010111010",
      "0100100001111110101011" when "0010111011",
      "0100100011011110101010" when "0010111100",
      "0100100100111110101010" when "0010111101",
      "0100100110011110101001" when "0010111110",
      "0100100111111110101000" when "0010111111",
      "0100101001011110100111" when "0011000000",
      "0100101010111110100110" when "0011000001",
      "0100101100011110100101" when "0011000010",
      "0100101101111110100100" when "0011000011",
      "0100101111011110100011" when "0011000100",
      "0100110000111110100010" when "0011000101",
      "0100110010011110100001" when "0011000110",
      "0100110011111110100000" when "0011000111",
      "0100110101011110011111" when "0011001000",
      "0100110110111110011110" when "0011001001",
      "0100111000011110011110" when "0011001010",
      "0100111001111110011101" when "0011001011",
      "0100111011011110011100" when "0011001100",
      "0100111100111110011011" when "0011001101",
      "0100111110011110011010" when "0011001110",
      "0100111111111110011001" when "0011001111",
      "0101000001011110011000" when "0011010000",
      "0101000010111110010111" when "0011010001",
      "0101000100011110010110" when "0011010010",
      "0101000101111110010101" when "0011010011",
      "0101000111011110010100" when "0011010100",
      "0101001000111110010011" when "0011010101",
      "0101001010011110010010" when "0011010110",
      "0101001011111110010001" when "0011010111",
      "0101001101011110010000" when "0011011000",
      "0101001110111110001111" when "0011011001",
      "0101010000011110001110" when "0011011010",
      "0101010001111110001101" when "0011011011",
      "0101010011011110001100" when "0011011100",
      "0101010100111110001010" when "0011011101",
      "0101010110011110001001" when "0011011110",
      "0101010111111110001000" when "0011011111",
      "0101011001011110000111" when "0011100000",
      "0101011010111110000110" when "0011100001",
      "0101011100011110000101" when "0011100010",
      "0101011101011110000100" when "0011100011",
      "0101011110111110000011" when "0011100100",
      "0101100000011110000010" when "0011100101",
      "0101100001111110000001" when "0011100110",
      "0101100011011110000000" when "0011100111",
      "0101100100111101111111" when "0011101000",
      "0101100110011101111110" when "0011101001",
      "0101100111111101111101" when "0011101010",
      "0101101001011101111011" when "0011101011",
      "0101101010111101111010" when "0011101100",
      "0101101100011101111001" when "0011101101",
      "0101101101111101111000" when "0011101110",
      "0101101111011101110111" when "0011101111",
      "0101110000111101110110" when "0011110000",
      "0101110010011101110101" when "0011110001",
      "0101110011111101110100" when "0011110010",
      "0101110100111101110010" when "0011110011",
      "0101110110011101110001" when "0011110100",
      "0101110111111101110000" when "0011110101",
      "0101111001011101101111" when "0011110110",
      "0101111010111101101110" when "0011110111",
      "0101111100011101101101" when "0011111000",
      "0101111101111101101011" when "0011111001",
      "0101111111011101101010" when "0011111010",
      "0110000000111101101001" when "0011111011",
      "0110000010011101101000" when "0011111100",
      "0110000011111101100111" when "0011111101",
      "0110000101011101100110" when "0011111110",
      "0110000110011101100100" when "0011111111",
      "0110000111111101100011" when "0100000000",
      "0110001001011101100010" when "0100000001",
      "0110001010111101100001" when "0100000010",
      "0110001100011101100000" when "0100000011",
      "0110001101111101011110" when "0100000100",
      "0110001111011101011101" when "0100000101",
      "0110010000111101011100" when "0100000110",
      "0110010010011101011011" when "0100000111",
      "0110010011111101011001" when "0100001000",
      "0110010100111101011000" when "0100001001",
      "0110010110011101010111" when "0100001010",
      "0110010111111101010110" when "0100001011",
      "0110011001011101010100" when "0100001100",
      "0110011010111101010011" when "0100001101",
      "0110011100011101010010" when "0100001110",
      "0110011101111101010001" when "0100001111",
      "0110011111011101001111" when "0100010000",
      "0110100000011101001110" when "0100010001",
      "0110100001111101001101" when "0100010010",
      "0110100011011101001100" when "0100010011",
      "0110100100111101001010" when "0100010100",
      "0110100110011101001001" when "0100010101",
      "0110100111111101001000" when "0100010110",
      "0110101001011101000110" when "0100010111",
      "0110101010011101000101" when "0100011000",
      "0110101011111101000100" when "0100011001",
      "0110101101011101000010" when "0100011010",
      "0110101110111101000001" when "0100011011",
      "0110110000011101000000" when "0100011100",
      "0110110001111100111110" when "0100011101",
      "0110110011011100111101" when "0100011110",
      "0110110100011100111100" when "0100011111",
      "0110110101111100111010" when "0100100000",
      "0110110111011100111001" when "0100100001",
      "0110111000111100111000" when "0100100010",
      "0110111010011100110110" when "0100100011",
      "0110111011111100110101" when "0100100100",
      "0110111100111100110100" when "0100100101",
      "0110111110011100110010" when "0100100110",
      "0110111111111100110001" when "0100100111",
      "0111000001011100110000" when "0100101000",
      "0111000010111100101110" when "0100101001",
      "0111000011111100101101" when "0100101010",
      "0111000101011100101011" when "0100101011",
      "0111000110111100101010" when "0100101100",
      "0111001000011100101001" when "0100101101",
      "0111001001111100100111" when "0100101110",
      "0111001011011100100110" when "0100101111",
      "0111001100011100100100" when "0100110000",
      "0111001101111100100011" when "0100110001",
      "0111001111011100100010" when "0100110010",
      "0111010000111100100000" when "0100110011",
      "0111010010011100011111" when "0100110100",
      "0111010011011100011101" when "0100110101",
      "0111010100111100011100" when "0100110110",
      "0111010110011100011010" when "0100110111",
      "0111010111111100011001" when "0100111000",
      "0111011001011100011000" when "0100111001",
      "0111011010011100010110" when "0100111010",
      "0111011011111100010101" when "0100111011",
      "0111011101011100010011" when "0100111100",
      "0111011110111100010010" when "0100111101",
      "0111011111111100010000" when "0100111110",
      "0111100001011100001111" when "0100111111",
      "0111100010111100001101" when "0101000000",
      "0111100100011100001100" when "0101000001",
      "0111100101011100001010" when "0101000010",
      "0111100110111100001001" when "0101000011",
      "0111101000011100000111" when "0101000100",
      "0111101001111100000110" when "0101000101",
      "0111101011011100000100" when "0101000110",
      "0111101100011100000011" when "0101000111",
      "0111101101111100000001" when "0101001000",
      "0111101111011100000000" when "0101001001",
      "0111110000111011111110" when "0101001010",
      "0111110001111011111101" when "0101001011",
      "0111110011011011111011" when "0101001100",
      "0111110100111011111010" when "0101001101",
      "0111110101111011111000" when "0101001110",
      "0111110111011011110111" when "0101001111",
      "0111111000111011110101" when "0101010000",
      "0111111010011011110100" when "0101010001",
      "0111111011011011110010" when "0101010010",
      "0111111100111011110000" when "0101010011",
      "0111111110011011101111" when "0101010100",
      "0111111111111011101101" when "0101010101",
      "1000000000111011101100" when "0101010110",
      "1000000010011011101010" when "0101010111",
      "1000000011111011101001" when "0101011000",
      "1000000100111011100111" when "0101011001",
      "1000000110011011100101" when "0101011010",
      "1000000111111011100100" when "0101011011",
      "1000001001011011100010" when "0101011100",
      "1000001010011011100001" when "0101011101",
      "1000001011111011011111" when "0101011110",
      "1000001101011011011101" when "0101011111",
      "1000001110011011011100" when "0101100000",
      "1000001111111011011010" when "0101100001",
      "1000010001011011011001" when "0101100010",
      "1000010010011011010111" when "0101100011",
      "1000010011111011010101" when "0101100100",
      "1000010101011011010100" when "0101100101",
      "1000010110011011010010" when "0101100110",
      "1000010111111011010000" when "0101100111",
      "1000011001011011001111" when "0101101000",
      "1000011010111011001101" when "0101101001",
      "1000011011111011001011" when "0101101010",
      "1000011101011011001010" when "0101101011",
      "1000011110111011001000" when "0101101100",
      "1000011111111011000110" when "0101101101",
      "1000100001011011000101" when "0101101110",
      "1000100010011011000011" when "0101101111",
      "1000100011111011000001" when "0101110000",
      "1000100101011011000000" when "0101110001",
      "1000100110011010111110" when "0101110010",
      "1000100111111010111100" when "0101110011",
      "1000101001011010111011" when "0101110100",
      "1000101010011010111001" when "0101110101",
      "1000101011111010110111" when "0101110110",
      "1000101101011010110110" when "0101110111",
      "1000101110011010110100" when "0101111000",
      "1000101111111010110010" when "0101111001",
      "1000110001011010110000" when "0101111010",
      "1000110010011010101111" when "0101111011",
      "1000110011111010101101" when "0101111100",
      "1000110100111010101011" when "0101111101",
      "1000110110011010101001" when "0101111110",
      "1000110111111010101000" when "0101111111",
      "1000111000111010100110" when "0110000000",
      "1000111010011010100100" when "0110000001",
      "1000111011011010100011" when "0110000010",
      "1000111100111010100001" when "0110000011",
      "1000111110011010011111" when "0110000100",
      "1000111111011010011101" when "0110000101",
      "1001000000111010011011" when "0110000110",
      "1001000001111010011010" when "0110000111",
      "1001000011011010011000" when "0110001000",
      "1001000100111010010110" when "0110001001",
      "1001000101111010010100" when "0110001010",
      "1001000111011010010011" when "0110001011",
      "1001001000011010010001" when "0110001100",
      "1001001001111010001111" when "0110001101",
      "1001001011011010001101" when "0110001110",
      "1001001100011010001011" when "0110001111",
      "1001001101111010001010" when "0110010000",
      "1001001110111010001000" when "0110010001",
      "1001010000011010000110" when "0110010010",
      "1001010001011010000100" when "0110010011",
      "1001010010111010000010" when "0110010100",
      "1001010011111010000001" when "0110010101",
      "1001010101011001111111" when "0110010110",
      "1001010110111001111101" when "0110010111",
      "1001010111111001111011" when "0110011000",
      "1001011001011001111001" when "0110011001",
      "1001011010011001110111" when "0110011010",
      "1001011011111001110101" when "0110011011",
      "1001011100111001110100" when "0110011100",
      "1001011110011001110010" when "0110011101",
      "1001011111011001110000" when "0110011110",
      "1001100000111001101110" when "0110011111",
      "1001100001111001101100" when "0110100000",
      "1001100011011001101010" when "0110100001",
      "1001100100011001101000" when "0110100010",
      "1001100101111001100111" when "0110100011",
      "1001100110111001100101" when "0110100100",
      "1001101000011001100011" when "0110100101",
      "1001101001011001100001" when "0110100110",
      "1001101010111001011111" when "0110100111",
      "1001101011111001011101" when "0110101000",
      "1001101101011001011011" when "0110101001",
      "1001101110011001011001" when "0110101010",
      "1001101111111001010111" when "0110101011",
      "1001110000111001010101" when "0110101100",
      "1001110010011001010100" when "0110101101",
      "1001110011011001010010" when "0110101110",
      "1001110100111001010000" when "0110101111",
      "1001110101111001001110" when "0110110000",
      "1001110111011001001100" when "0110110001",
      "1001111000011001001010" when "0110110010",
      "1001111001111001001000" when "0110110011",
      "1001111010111001000110" when "0110110100",
      "1001111100011001000100" when "0110110101",
      "1001111101011001000010" when "0110110110",
      "1001111110111001000000" when "0110110111",
      "1001111111111000111110" when "0110111000",
      "1010000001011000111100" when "0110111001",
      "1010000010011000111010" when "0110111010",
      "1010000011011000111000" when "0110111011",
      "1010000100111000110110" when "0110111100",
      "1010000101111000110100" when "0110111101",
      "1010000111011000110010" when "0110111110",
      "1010001000011000110000" when "0110111111",
      "1010001001111000101110" when "0111000000",
      "1010001010111000101100" when "0111000001",
      "1010001011111000101010" when "0111000010",
      "1010001101011000101000" when "0111000011",
      "1010001110011000100110" when "0111000100",
      "1010001111111000100100" when "0111000101",
      "1010010000111000100010" when "0111000110",
      "1010010010011000100000" when "0111000111",
      "1010010011011000011110" when "0111001000",
      "1010010100011000011100" when "0111001001",
      "1010010101111000011010" when "0111001010",
      "1010010110111000011000" when "0111001011",
      "1010011000011000010110" when "0111001100",
      "1010011001011000010100" when "0111001101",
      "1010011010011000010010" when "0111001110",
      "1010011011111000010000" when "0111001111",
      "1010011100111000001110" when "0111010000",
      "1010011101111000001100" when "0111010001",
      "1010011111011000001010" when "0111010010",
      "1010100000011000001000" when "0111010011",
      "1010100001111000000110" when "0111010100",
      "1010100010111000000100" when "0111010101",
      "1010100011111000000010" when "0111010110",
      "1010100101011000000000" when "0111010111",
      "1010100110010111111101" when "0111011000",
      "1010100111010111111011" when "0111011001",
      "1010101000110111111001" when "0111011010",
      "1010101001110111110111" when "0111011011",
      "1010101010110111110101" when "0111011100",
      "1010101100010111110011" when "0111011101",
      "1010101101010111110001" when "0111011110",
      "1010101110010111101111" when "0111011111",
      "1010101111110111101101" when "0111100000",
      "1010110000110111101011" when "0111100001",
      "1010110001110111101001" when "0111100010",
      "1010110011010111100110" when "0111100011",
      "1010110100010111100100" when "0111100100",
      "1010110101010111100010" when "0111100101",
      "1010110110110111100000" when "0111100110",
      "1010110111110111011110" when "0111100111",
      "1010111000110111011100" when "0111101000",
      "1010111001110111011010" when "0111101001",
      "1010111011010111010111" when "0111101010",
      "1010111100010111010101" when "0111101011",
      "1010111101010111010011" when "0111101100",
      "1010111110110111010001" when "0111101101",
      "1010111111110111001111" when "0111101110",
      "1011000000110111001101" when "0111101111",
      "1011000001110111001011" when "0111110000",
      "1011000011010111001000" when "0111110001",
      "1011000100010111000110" when "0111110010",
      "1011000101010111000100" when "0111110011",
      "1011000110110111000010" when "0111110100",
      "1011000111110111000000" when "0111110101",
      "1011001000110110111101" when "0111110110",
      "1011001001110110111011" when "0111110111",
      "1011001011010110111001" when "0111111000",
      "1011001100010110110111" when "0111111001",
      "1011001101010110110101" when "0111111010",
      "1011001110010110110011" when "0111111011",
      "1011001111110110110000" when "0111111100",
      "1011010000110110101110" when "0111111101",
      "1011010001110110101100" when "0111111110",
      "1011010010110110101010" when "0111111111",
      "1011010011110110100111" when "1000000000",
      "1011010101010110100101" when "1000000001",
      "1011010110010110100011" when "1000000010",
      "1011010111010110100001" when "1000000011",
      "1011011000010110011111" when "1000000100",
      "1011011001110110011100" when "1000000101",
      "1011011010110110011010" when "1000000110",
      "1011011011110110011000" when "1000000111",
      "1011011100110110010110" when "1000001000",
      "1011011101110110010011" when "1000001001",
      "1011011110110110010001" when "1000001010",
      "1011100000010110001111" when "1000001011",
      "1011100001010110001101" when "1000001100",
      "1011100010010110001010" when "1000001101",
      "1011100011010110001000" when "1000001110",
      "1011100100010110000110" when "1000001111",
      "1011100101110110000011" when "1000010000",
      "1011100110110110000001" when "1000010001",
      "1011100111110101111111" when "1000010010",
      "1011101000110101111101" when "1000010011",
      "1011101001110101111010" when "1000010100",
      "1011101010110101111000" when "1000010101",
      "1011101011110101110110" when "1000010110",
      "1011101101010101110011" when "1000010111",
      "1011101110010101110001" when "1000011000",
      "1011101111010101101111" when "1000011001",
      "1011110000010101101101" when "1000011010",
      "1011110001010101101010" when "1000011011",
      "1011110010010101101000" when "1000011100",
      "1011110011010101100110" when "1000011101",
      "1011110100110101100011" when "1000011110",
      "1011110101110101100001" when "1000011111",
      "1011110110110101011111" when "1000100000",
      "1011110111110101011100" when "1000100001",
      "1011111000110101011010" when "1000100010",
      "1011111001110101011000" when "1000100011",
      "1011111010110101010101" when "1000100100",
      "1011111011110101010011" when "1000100101",
      "1011111100110101010001" when "1000100110",
      "1011111101110101001110" when "1000100111",
      "1011111110110101001100" when "1000101000",
      "1100000000010101001010" when "1000101001",
      "1100000001010101000111" when "1000101010",
      "1100000010010101000101" when "1000101011",
      "1100000011010101000011" when "1000101100",
      "1100000100010101000000" when "1000101101",
      "1100000101010100111110" when "1000101110",
      "1100000110010100111011" when "1000101111",
      "1100000111010100111001" when "1000110000",
      "1100001000010100110111" when "1000110001",
      "1100001001010100110100" when "1000110010",
      "1100001010010100110010" when "1000110011",
      "1100001011010100110000" when "1000110100",
      "1100001100010100101101" when "1000110101",
      "1100001101010100101011" when "1000110110",
      "1100001110010100101000" when "1000110111",
      "1100001111010100100110" when "1000111000",
      "1100010000010100100100" when "1000111001",
      "1100010001010100100001" when "1000111010",
      "1100010010010100011111" when "1000111011",
      "1100010011010100011100" when "1000111100",
      "1100010100010100011010" when "1000111101",
      "1100010101010100010111" when "1000111110",
      "1100010110010100010101" when "1000111111",
      "1100010111010100010011" when "1001000000",
      "1100011000010100010000" when "1001000001",
      "1100011001010100001110" when "1001000010",
      "1100011010010100001011" when "1001000011",
      "1100011011010100001001" when "1001000100",
      "1100011100010100000110" when "1001000101",
      "1100011101010100000100" when "1001000110",
      "1100011110010100000010" when "1001000111",
      "1100011111010011111111" when "1001001000",
      "1100100000010011111101" when "1001001001",
      "1100100001010011111010" when "1001001010",
      "1100100010010011111000" when "1001001011",
      "1100100011010011110101" when "1001001100",
      "1100100100010011110011" when "1001001101",
      "1100100101010011110000" when "1001001110",
      "1100100110010011101110" when "1001001111",
      "1100100111010011101011" when "1001010000",
      "1100101000010011101001" when "1001010001",
      "1100101001010011100110" when "1001010010",
      "1100101010010011100100" when "1001010011",
      "1100101010110011100001" when "1001010100",
      "1100101011110011011111" when "1001010101",
      "1100101100110011011100" when "1001010110",
      "1100101101110011011010" when "1001010111",
      "1100101110110011010111" when "1001011000",
      "1100101111110011010101" when "1001011001",
      "1100110000110011010010" when "1001011010",
      "1100110001110011010000" when "1001011011",
      "1100110010110011001101" when "1001011100",
      "1100110011110011001011" when "1001011101",
      "1100110100010011001000" when "1001011110",
      "1100110101010011000110" when "1001011111",
      "1100110110010011000011" when "1001100000",
      "1100110111010011000001" when "1001100001",
      "1100111000010010111110" when "1001100010",
      "1100111001010010111100" when "1001100011",
      "1100111010010010111001" when "1001100100",
      "1100111010110010110111" when "1001100101",
      "1100111011110010110100" when "1001100110",
      "1100111100110010110010" when "1001100111",
      "1100111101110010101111" when "1001101000",
      "1100111110110010101101" when "1001101001",
      "1100111111110010101010" when "1001101010",
      "1101000000110010100111" when "1001101011",
      "1101000001010010100101" when "1001101100",
      "1101000010010010100010" when "1001101101",
      "1101000011010010100000" when "1001101110",
      "1101000100010010011101" when "1001101111",
      "1101000101010010011011" when "1001110000",
      "1101000101110010011000" when "1001110001",
      "1101000110110010010110" when "1001110010",
      "1101000111110010010011" when "1001110011",
      "1101001000110010010000" when "1001110100",
      "1101001001110010001110" when "1001110101",
      "1101001010010010001011" when "1001110110",
      "1101001011010010001001" when "1001110111",
      "1101001100010010000110" when "1001111000",
      "1101001101010010000011" when "1001111001",
      "1101001101110010000001" when "1001111010",
      "1101001110110001111110" when "1001111011",
      "1101001111110001111100" when "1001111100",
      "1101010000110001111001" when "1001111101",
      "1101010001110001110110" when "1001111110",
      "1101010010010001110100" when "1001111111",
      "1101010011010001110001" when "1010000000",
      "1101010100010001101111" when "1010000001",
      "1101010100110001101100" when "1010000010",
      "1101010101110001101001" when "1010000011",
      "1101010110110001100111" when "1010000100",
      "1101010111110001100100" when "1010000101",
      "1101011000010001100010" when "1010000110",
      "1101011001010001011111" when "1010000111",
      "1101011010010001011100" when "1010001000",
      "1101011011010001011010" when "1010001001",
      "1101011011110001010111" when "1010001010",
      "1101011100110001010100" when "1010001011",
      "1101011101110001010010" when "1010001100",
      "1101011110010001001111" when "1010001101",
      "1101011111010001001100" when "1010001110",
      "1101100000010001001010" when "1010001111",
      "1101100000110001000111" when "1010010000",
      "1101100001110001000100" when "1010010001",
      "1101100010110001000010" when "1010010010",
      "1101100011010000111111" when "1010010011",
      "1101100100010000111101" when "1010010100",
      "1101100101010000111010" when "1010010101",
      "1101100101110000110111" when "1010010110",
      "1101100110110000110101" when "1010010111",
      "1101100111110000110010" when "1010011000",
      "1101101000010000101111" when "1010011001",
      "1101101001010000101100" when "1010011010",
      "1101101010010000101010" when "1010011011",
      "1101101010110000100111" when "1010011100",
      "1101101011110000100100" when "1010011101",
      "1101101100110000100010" when "1010011110",
      "1101101101010000011111" when "1010011111",
      "1101101110010000011100" when "1010100000",
      "1101101110110000011010" when "1010100001",
      "1101101111110000010111" when "1010100010",
      "1101110000110000010100" when "1010100011",
      "1101110001010000010010" when "1010100100",
      "1101110010010000001111" when "1010100101",
      "1101110010110000001100" when "1010100110",
      "1101110011110000001001" when "1010100111",
      "1101110100110000000111" when "1010101000",
      "1101110101010000000100" when "1010101001",
      "1101110110010000000001" when "1010101010",
      "1101110110101111111111" when "1010101011",
      "1101110111101111111100" when "1010101100",
      "1101111000001111111001" when "1010101101",
      "1101111001001111110110" when "1010101110",
      "1101111010001111110100" when "1010101111",
      "1101111010101111110001" when "1010110000",
      "1101111011101111101110" when "1010110001",
      "1101111100001111101011" when "1010110010",
      "1101111101001111101001" when "1010110011",
      "1101111101101111100110" when "1010110100",
      "1101111110101111100011" when "1010110101",
      "1101111111001111100001" when "1010110110",
      "1110000000001111011110" when "1010110111",
      "1110000000101111011011" when "1010111000",
      "1110000001101111011000" when "1010111001",
      "1110000010001111010110" when "1010111010",
      "1110000011001111010011" when "1010111011",
      "1110000011101111010000" when "1010111100",
      "1110000100101111001101" when "1010111101",
      "1110000101001111001010" when "1010111110",
      "1110000110001111001000" when "1010111111",
      "1110000110101111000101" when "1011000000",
      "1110000111101111000010" when "1011000001",
      "1110001000001110111111" when "1011000010",
      "1110001001001110111101" when "1011000011",
      "1110001001101110111010" when "1011000100",
      "1110001010101110110111" when "1011000101",
      "1110001011001110110100" when "1011000110",
      "1110001100001110110010" when "1011000111",
      "1110001100101110101111" when "1011001000",
      "1110001101001110101100" when "1011001001",
      "1110001110001110101001" when "1011001010",
      "1110001110101110100110" when "1011001011",
      "1110001111101110100100" when "1011001100",
      "1110010000001110100001" when "1011001101",
      "1110010001001110011110" when "1011001110",
      "1110010001101110011011" when "1011001111",
      "1110010010001110011000" when "1011010000",
      "1110010011001110010110" when "1011010001",
      "1110010011101110010011" when "1011010010",
      "1110010100101110010000" when "1011010011",
      "1110010101001110001101" when "1011010100",
      "1110010101101110001010" when "1011010101",
      "1110010110101110000111" when "1011010110",
      "1110010111001110000101" when "1011010111",
      "1110011000001110000010" when "1011011000",
      "1110011000101101111111" when "1011011001",
      "1110011001001101111100" when "1011011010",
      "1110011010001101111001" when "1011011011",
      "1110011010101101110111" when "1011011100",
      "1110011011001101110100" when "1011011101",
      "1110011100001101110001" when "1011011110",
      "1110011100101101101110" when "1011011111",
      "1110011101001101101011" when "1011100000",
      "1110011110001101101000" when "1011100001",
      "1110011110101101100110" when "1011100010",
      "1110011111001101100011" when "1011100011",
      "1110100000001101100000" when "1011100100",
      "1110100000101101011101" when "1011100101",
      "1110100001001101011010" when "1011100110",
      "1110100010001101010111" when "1011100111",
      "1110100010101101010100" when "1011101000",
      "1110100011001101010010" when "1011101001",
      "1110100100001101001111" when "1011101010",
      "1110100100101101001100" when "1011101011",
      "1110100101001101001001" when "1011101100",
      "1110100110001101000110" when "1011101101",
      "1110100110101101000011" when "1011101110",
      "1110100111001101000000" when "1011101111",
      "1110100111101100111110" when "1011110000",
      "1110101000101100111011" when "1011110001",
      "1110101001001100111000" when "1011110010",
      "1110101001101100110101" when "1011110011",
      "1110101010001100110010" when "1011110100",
      "1110101011001100101111" when "1011110101",
      "1110101011101100101100" when "1011110110",
      "1110101100001100101001" when "1011110111",
      "1110101100101100100111" when "1011111000",
      "1110101101101100100100" when "1011111001",
      "1110101110001100100001" when "1011111010",
      "1110101110101100011110" when "1011111011",
      "1110101111001100011011" when "1011111100",
      "1110110000001100011000" when "1011111101",
      "1110110000101100010101" when "1011111110",
      "1110110001001100010010" when "1011111111",
      "1110110001101100001111" when "1100000000",
      "1110110010001100001100" when "1100000001",
      "1110110011001100001010" when "1100000010",
      "1110110011101100000111" when "1100000011",
      "1110110100001100000100" when "1100000100",
      "1110110100101100000001" when "1100000101",
      "1110110101001011111110" when "1100000110",
      "1110110101101011111011" when "1100000111",
      "1110110110101011111000" when "1100001000",
      "1110110111001011110101" when "1100001001",
      "1110110111101011110010" when "1100001010",
      "1110111000001011101111" when "1100001011",
      "1110111000101011101100" when "1100001100",
      "1110111001001011101001" when "1100001101",
      "1110111010001011100111" when "1100001110",
      "1110111010101011100100" when "1100001111",
      "1110111011001011100001" when "1100010000",
      "1110111011101011011110" when "1100010001",
      "1110111100001011011011" when "1100010010",
      "1110111100101011011000" when "1100010011",
      "1110111101001011010101" when "1100010100",
      "1110111101101011010010" when "1100010101",
      "1110111110101011001111" when "1100010110",
      "1110111111001011001100" when "1100010111",
      "1110111111101011001001" when "1100011000",
      "1111000000001011000110" when "1100011001",
      "1111000000101011000011" when "1100011010",
      "1111000001001011000000" when "1100011011",
      "1111000001101010111101" when "1100011100",
      "1111000010001010111010" when "1100011101",
      "1111000010101010111000" when "1100011110",
      "1111000011001010110101" when "1100011111",
      "1111000011101010110010" when "1100100000",
      "1111000100001010101111" when "1100100001",
      "1111000100101010101100" when "1100100010",
      "1111000101001010101001" when "1100100011",
      "1111000110001010100110" when "1100100100",
      "1111000110101010100011" when "1100100101",
      "1111000111001010100000" when "1100100110",
      "1111000111101010011101" when "1100100111",
      "1111001000001010011010" when "1100101000",
      "1111001000101010010111" when "1100101001",
      "1111001001001010010100" when "1100101010",
      "1111001001101010010001" when "1100101011",
      "1111001010001010001110" when "1100101100",
      "1111001010101010001011" when "1100101101",
      "1111001011001010001000" when "1100101110",
      "1111001011101010000101" when "1100101111",
      "1111001100001010000010" when "1100110000",
      "1111001100101001111111" when "1100110001",
      "1111001101001001111100" when "1100110010",
      "1111001101101001111001" when "1100110011",
      "1111001110001001110110" when "1100110100",
      "1111001110101001110011" when "1100110101",
      "1111001111001001110000" when "1100110110",
      "1111001111001001101101" when "1100110111",
      "1111001111101001101010" when "1100111000",
      "1111010000001001100111" when "1100111001",
      "1111010000101001100100" when "1100111010",
      "1111010001001001100001" when "1100111011",
      "1111010001101001011110" when "1100111100",
      "1111010010001001011011" when "1100111101",
      "1111010010101001011000" when "1100111110",
      "1111010011001001010101" when "1100111111",
      "1111010011101001010010" when "1101000000",
      "1111010100001001001111" when "1101000001",
      "1111010100101001001100" when "1101000010",
      "1111010101001001001001" when "1101000011",
      "1111010101001001000110" when "1101000100",
      "1111010101101001000011" when "1101000101",
      "1111010110001001000000" when "1101000110",
      "1111010110101000111101" when "1101000111",
      "1111010111001000111010" when "1101001000",
      "1111010111101000110111" when "1101001001",
      "1111011000001000110100" when "1101001010",
      "1111011000101000110001" when "1101001011",
      "1111011000101000101110" when "1101001100",
      "1111011001001000101011" when "1101001101",
      "1111011001101000101000" when "1101001110",
      "1111011010001000100101" when "1101001111",
      "1111011010101000100010" when "1101010000",
      "1111011011001000011111" when "1101010001",
      "1111011011101000011100" when "1101010010",
      "1111011011101000011001" when "1101010011",
      "1111011100001000010110" when "1101010100",
      "1111011100101000010011" when "1101010101",
      "1111011101001000010000" when "1101010110",
      "1111011101101000001101" when "1101010111",
      "1111011101101000001010" when "1101011000",
      "1111011110001000000111" when "1101011001",
      "1111011110101000000100" when "1101011010",
      "1111011111001000000001" when "1101011011",
      "1111011111100111111110" when "1101011100",
      "1111011111100111111011" when "1101011101",
      "1111100000000111110111" when "1101011110",
      "1111100000100111110100" when "1101011111",
      "1111100001000111110001" when "1101100000",
      "1111100001000111101110" when "1101100001",
      "1111100001100111101011" when "1101100010",
      "1111100010000111101000" when "1101100011",
      "1111100010100111100101" when "1101100100",
      "1111100010100111100010" when "1101100101",
      "1111100011000111011111" when "1101100110",
      "1111100011100111011100" when "1101100111",
      "1111100100000111011001" when "1101101000",
      "1111100100000111010110" when "1101101001",
      "1111100100100111010011" when "1101101010",
      "1111100101000111010000" when "1101101011",
      "1111100101000111001101" when "1101101100",
      "1111100101100111001010" when "1101101101",
      "1111100110000111000111" when "1101101110",
      "1111100110100111000100" when "1101101111",
      "1111100110100111000001" when "1101110000",
      "1111100111000110111101" when "1101110001",
      "1111100111100110111010" when "1101110010",
      "1111100111100110110111" when "1101110011",
      "1111101000000110110100" when "1101110100",
      "1111101000100110110001" when "1101110101",
      "1111101000100110101110" when "1101110110",
      "1111101001000110101011" when "1101110111",
      "1111101001100110101000" when "1101111000",
      "1111101001100110100101" when "1101111001",
      "1111101010000110100010" when "1101111010",
      "1111101010100110011111" when "1101111011",
      "1111101010100110011100" when "1101111100",
      "1111101011000110011001" when "1101111101",
      "1111101011000110010110" when "1101111110",
      "1111101011100110010010" when "1101111111",
      "1111101100000110001111" when "1110000000",
      "1111101100000110001100" when "1110000001",
      "1111101100100110001001" when "1110000010",
      "1111101100100110000110" when "1110000011",
      "1111101101000110000011" when "1110000100",
      "1111101101100110000000" when "1110000101",
      "1111101101100101111101" when "1110000110",
      "1111101110000101111010" when "1110000111",
      "1111101110000101110111" when "1110001000",
      "1111101110100101110100" when "1110001001",
      "1111101111000101110001" when "1110001010",
      "1111101111000101101101" when "1110001011",
      "1111101111100101101010" when "1110001100",
      "1111101111100101100111" when "1110001101",
      "1111110000000101100100" when "1110001110",
      "1111110000000101100001" when "1110001111",
      "1111110000100101011110" when "1110010000",
      "1111110000100101011011" when "1110010001",
      "1111110001000101011000" when "1110010010",
      "1111110001000101010101" when "1110010011",
      "1111110001100101010010" when "1110010100",
      "1111110001100101001110" when "1110010101",
      "1111110010000101001011" when "1110010110",
      "1111110010100101001000" when "1110010111",
      "1111110010100101000101" when "1110011000",
      "1111110011000101000010" when "1110011001",
      "1111110011000100111111" when "1110011010",
      "1111110011000100111100" when "1110011011",
      "1111110011100100111001" when "1110011100",
      "1111110011100100110110" when "1110011101",
      "1111110100000100110011" when "1110011110",
      "1111110100000100101111" when "1110011111",
      "1111110100100100101100" when "1110100000",
      "1111110100100100101001" when "1110100001",
      "1111110101000100100110" when "1110100010",
      "1111110101000100100011" when "1110100011",
      "1111110101100100100000" when "1110100100",
      "1111110101100100011101" when "1110100101",
      "1111110110000100011010" when "1110100110",
      "1111110110000100010111" when "1110100111",
      "1111110110000100010011" when "1110101000",
      "1111110110100100010000" when "1110101001",
      "1111110110100100001101" when "1110101010",
      "1111110111000100001010" when "1110101011",
      "1111110111000100000111" when "1110101100",
      "1111110111000100000100" when "1110101101",
      "1111110111100100000001" when "1110101110",
      "1111110111100011111110" when "1110101111",
      "1111111000000011111011" when "1110110000",
      "1111111000000011110111" when "1110110001",
      "1111111000000011110100" when "1110110010",
      "1111111000100011110001" when "1110110011",
      "1111111000100011101110" when "1110110100",
      "1111111000100011101011" when "1110110101",
      "1111111001000011101000" when "1110110110",
      "1111111001000011100101" when "1110110111",
      "1111111001100011100010" when "1110111000",
      "1111111001100011011111" when "1110111001",
      "1111111001100011011011" when "1110111010",
      "1111111010000011011000" when "1110111011",
      "1111111010000011010101" when "1110111100",
      "1111111010000011010010" when "1110111101",
      "1111111010100011001111" when "1110111110",
      "1111111010100011001100" when "1110111111",
      "1111111010100011001001" when "1111000000",
      "1111111010100011000110" when "1111000001",
      "1111111011000011000010" when "1111000010",
      "1111111011000010111111" when "1111000011",
      "1111111011000010111100" when "1111000100",
      "1111111011100010111001" when "1111000101",
      "1111111011100010110110" when "1111000110",
      "1111111011100010110011" when "1111000111",
      "1111111011100010110000" when "1111001000",
      "1111111100000010101100" when "1111001001",
      "1111111100000010101001" when "1111001010",
      "1111111100000010100110" when "1111001011",
      "1111111100000010100011" when "1111001100",
      "1111111100100010100000" when "1111001101",
      "1111111100100010011101" when "1111001110",
      "1111111100100010011010" when "1111001111",
      "1111111100100010010111" when "1111010000",
      "1111111101000010010011" when "1111010001",
      "1111111101000010010000" when "1111010010",
      "1111111101000010001101" when "1111010011",
      "1111111101000010001010" when "1111010100",
      "1111111101100010000111" when "1111010101",
      "1111111101100010000100" when "1111010110",
      "1111111101100010000001" when "1111010111",
      "1111111101100001111110" when "1111011000",
      "1111111101100001111010" when "1111011001",
      "1111111110000001110111" when "1111011010",
      "1111111110000001110100" when "1111011011",
      "1111111110000001110001" when "1111011100",
      "1111111110000001101110" when "1111011101",
      "1111111110000001101011" when "1111011110",
      "1111111110000001101000" when "1111011111",
      "1111111110100001100100" when "1111100000",
      "1111111110100001100001" when "1111100001",
      "1111111110100001011110" when "1111100010",
      "1111111110100001011011" when "1111100011",
      "1111111110100001011000" when "1111100100",
      "1111111110100001010101" when "1111100101",
      "1111111110100001010010" when "1111100110",
      "1111111110100001001110" when "1111100111",
      "1111111111000001001011" when "1111101000",
      "1111111111000001001000" when "1111101001",
      "1111111111000001000101" when "1111101010",
      "1111111111000001000010" when "1111101011",
      "1111111111000000111111" when "1111101100",
      "1111111111000000111100" when "1111101101",
      "1111111111000000111001" when "1111101110",
      "1111111111000000110101" when "1111101111",
      "1111111111000000110010" when "1111110000",
      "1111111111000000101111" when "1111110001",
      "1111111111100000101100" when "1111110010",
      "1111111111100000101001" when "1111110011",
      "1111111111100000100110" when "1111110100",
      "1111111111100000100011" when "1111110101",
      "1111111111100000011111" when "1111110110",
      "1111111111100000011100" when "1111110111",
      "1111111111100000011001" when "1111111000",
      "1111111111100000010110" when "1111111001",
      "1111111111100000010011" when "1111111010",
      "1111111111100000010000" when "1111111011",
      "1111111111100000001101" when "1111111100",
      "1111111111100000001001" when "1111111101",
      "1111111111100000000110" when "1111111110",
      "1111111111100000000011" when "1111111111",
      "----------------------" when others;
   Y1 <= Y0_d1; -- for the possible blockram register
   Y <= Y1;
end architecture;

--------------------------------------------------------------------------------
--                                FixSinCos_11
--                    (FixSinCosPoly_LSBm11_Freq200_uid2)
-- VHDL generated for DummyFPGA @ 200MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Antoine Martinet, Guillaume Sergent, (2013-2019)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles
-- Clock period (ns): 5
-- Target frequency (MHz): 200
-- Input signals: X
-- Output signals: S C
--  approx. input signal timings: X: (c0, 0.000000ns)
--  approx. output signal timings: S: (c1, 2.239062ns)C: (c1, 2.239062ns)

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixSinCos_11 is
    port (clk, rst : in std_logic;
          X : in  std_logic_vector(11 downto 0);
          S : out  std_logic_vector(11 downto 0);
          C : out  std_logic_vector(11 downto 0)   );
end entity;

architecture arch of FixSinCos_11 is
   component SinCosTable_Freq200_uid4 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(9 downto 0);
             Y : out  std_logic_vector(21 downto 0)   );
   end component;

signal X_sgn, X_sgn_d1 :  std_logic;
   -- timing of X_sgn: (c0, 0.000000ns)
signal Q, Q_d1 :  std_logic;
   -- timing of Q: (c0, 0.000000ns)
signal sinCosTabIn :  std_logic_vector(9 downto 0);
   -- timing of sinCosTabIn: (c0, 0.000000ns)
signal C_sgn, C_sgn_d1 :  std_logic;
   -- timing of C_sgn: (c0, 0.000000ns)
signal SinCos :  std_logic_vector(21 downto 0);
   -- timing of SinCos: (c1, 2.239062ns)
signal S_out :  std_logic_vector(10 downto 0);
   -- timing of S_out: (c1, 2.239062ns)
signal C_out :  std_logic_vector(10 downto 0);
   -- timing of C_out: (c1, 2.239062ns)
signal S_wo_sgn :  std_logic_vector(10 downto 0);
   -- timing of S_wo_sgn: (c1, 2.239062ns)
signal C_wo_sgn :  std_logic_vector(10 downto 0);
   -- timing of C_wo_sgn: (c1, 2.239062ns)
signal S_wo_sgn_ext :  std_logic_vector(11 downto 0);
   -- timing of S_wo_sgn_ext: (c1, 2.239062ns)
signal C_wo_sgn_ext :  std_logic_vector(11 downto 0);
   -- timing of C_wo_sgn_ext: (c1, 2.239062ns)
signal S_wo_sgn_neg :  std_logic_vector(11 downto 0);
   -- timing of S_wo_sgn_neg: (c1, 2.239062ns)
signal C_wo_sgn_neg :  std_logic_vector(11 downto 0);
   -- timing of C_wo_sgn_neg: (c1, 2.239062ns)
begin
   process(clk, rst)
      begin
         if rst = '1' then
            X_sgn_d1 <=  '0';
            Q_d1 <=  '0';
            C_sgn_d1 <=  '0';
         elsif clk'event and clk = '1' then
            X_sgn_d1 <=  X_sgn;
            Q_d1 <=  Q;
            C_sgn_d1 <=  C_sgn;
         end if;
      end process;
   X_sgn <= X(11);
   Q <= X(10);
   sinCosTabIn <= X (9 downto 0);
   C_sgn <= Q xor X_sgn;
   SinCosTable: SinCosTable_Freq200_uid4
      port map ( clk  => clk,
                 rst  => rst,
                 X => sinCosTabIn,
                 Y => SinCos);
   S_out <= SinCos(21 downto 11);
   C_out <= SinCos(10 downto 0);
   S_wo_sgn <= C_out when Q_d1 = '1' else S_out;
   C_wo_sgn <= S_out when Q_d1 = '1' else C_out;
   S_wo_sgn_ext <= '0' & S_wo_sgn;
   C_wo_sgn_ext <= '0' & C_wo_sgn;
   S_wo_sgn_neg <= (not S_wo_sgn_ext) + 1;
   C_wo_sgn_neg <= (not C_wo_sgn_ext) + 1;
   S <= S_wo_sgn_ext when X_sgn_d1 = '0' else S_wo_sgn_neg;
   C <= C_wo_sgn_ext when C_sgn_d1 = '0' else C_wo_sgn_neg;
end architecture;

